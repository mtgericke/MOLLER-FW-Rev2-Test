-------------------------------------------------------------
-- Filename:  LFSR11PROM.VHD
-- Authors: 
-- 	from http://www.xilinx.com/support/documentation/sw_manuals/xilinx14_4/xst_v6s6.pdf  p262
--		Alain Zarembowitch / MSS
-- Version: Rev 0
-- Last modified: 8/24/16

-- Inheritance: 	ROM1.VHD
--
-- description:  synthesizable generic dual port ROM. Customized for LFSR11P.
-- Warning: convoluted pointers to alleviate re-writing the ROM contents transferred from a Xilinx block ram.
---------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity LFSR11PROM is
	 Generic (
		DATA_WIDTH: integer := 8;	
		ADDR_WIDTH: integer := 11
	);
    Port ( 
	    -- Port A
		CLKA   : in  std_logic;
		CSA: in std_logic;	-- chip select, active high
		OEA : in std_logic;	-- output enable, active high
		ADDRA  : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		DOA  : out std_logic_vector(DATA_WIDTH-1 downto 0);
			-- Stores 8 contiguous PRBS-11 sequence in DATA_OUT(7:0). Period is 8*2047 bits.	
			-- SOF is placed in DATA_OUT(8)

		-- Port B 
		CLKB   : in  std_logic;
		CSB: in std_logic;	-- chip select, active high
		OEB : in std_logic;	-- output enable, active high
		ADDRB  : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		DOB  : out std_logic_vector(DATA_WIDTH-1 downto 0)
		);
end entity;

architecture Behavioral of LFSR11PROM is
--------------------------------------------------------
--     SIGNALS
--------------------------------------------------------
-- inferred rom
signal DOA_local: std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
signal DOB_local: std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
type ROM_TYPE is array ( (2**(ADDR_WIDTH-5))-1 downto 0 ) of std_logic_vector(255 downto 0);
constant ROM : ROM_TYPE := (
      -- Address 0 to 511
      x"3BA0CC2D85C4380D2E8334476B74B90E82C970180CD3B4473F01CE7CF8F31F00",
      x"114F7EFC53B5BBA09858F2B64237419B0BDF54B8F3B5BA0872B6164236E971E5",
      x"EE7D05C46C7859F14E7D046C8696BD053AA33412B6E925904CD2B617EADC0795",
      x"15111B0B8B21CF81CF80676A898E7DFAA3CADDFAA2623714469643CA76E873B5",
      x"FD504D8493B5456FD413B5111AA361CF2B75BB5E5714B9F1E56FD5BB5FFFFE57",
      x"76E9DB5F0099F1B0B24827C131E5911AF714B8590F81314F2B21CE29256E839E",
      x"CE839F55BAA36067C19B5FAA23CA898FD5104D2E298E7C524924390ED6BC076A",
      x"66961617EB74ED7BF5BB0A2263CB8BDF00CD84C7C0321DAE29DA09253B5E0361",
      x"7740995B0A89711A5C06698ED6E8721D0493E13018A6698F7E029CF9F0E73F00",
      x"239EFCF8A76A774131B1E46D856E823617BEA970E76B7511E46C2D846CD2E3CA",
      x"DDFB0A88D9F0B2E29DFA08D80C2D7B0B744669246CD34B2099A46D2FD4B90F2A",
      X"2A22361616439E039F01CFD4121DFBF44795BBF545C56E288C2C8794EDD0E76A",
      X"FBA19A08276B8BDEA8276A233446C39E57EA76BDAE2872E3CBDFAA77BFFEFDAF",
      X"ECD2B7BF0032E36165914E8263CA2335EE2970B31E02639E56429C534ADC063D",
      X"9C073FAB7447C1CE8237BF544794131FAB219A5C521CF9A49248721CAC790FD4",
      X"CC2C2D2ED6E9DAF7EA771544C69617BF019A098F81653A5C53B4134A76BC06C2",
      -- Address 512 to 1023
      X"EF8032B71412E334B80CD21CADD1E53A0826C361304CD31EFD0438F3E1CF7F00",
      X"463CF9F14FD5EE826262C9DB0ADD046D2E7C53E1CED7EA22C8D95A08D9A4C795",
      X"BAF71510B3E165C53BF511B0195AF616E88CD248D8A697403249DB5EA8731F54",
      X"55446C2C2C863C073E039EA9253AF6E98F2A77EB8B8ADD5018590E29DBA1CFD5",
      X"F64335114ED616BD514FD446688C863DAFD4ED7A5D51E4C697BF55EF7EFDFB5F",
      X"D9A56F7F0164C6C3CA229D04C794476ADC53E0663D04C63CAD8438A794B80D7A",
      X"390F7E56E98E829D056F7EA98E28273E564334B9A438F2492591E43858F31EA8",
      X"98595A5CACD3B5EFD5EF2A888C2D2F7E0334131E03CB74B8A6682794EC780D84",
      X"DF01656E2924C6697019A4395AA3CB75104C86C36098A63DFA0970E6C39FFF00",
      X"8C78F2E39FAADD05C5C492B715BA09DA5CF8A6C29DAFD54590B3B510B2498F2B",
      X"75EF2B2066C3CB8A77EA236033B4EC2DD019A591B04D2F816492B6BD50E73EA8",
      X"AA88D858580C790E7C063C534B74ECD31F55EED61715BBA130B21C52B6439FAB",
      X"EC876A229CAC2D7AA39EA88DD0180D7B5EA9DBF5BAA2C88D2F7FABDEFDFAF7BF",
      X"B34BDFFE02C88C8795453A098E298FD4B8A7C0CD7A088C795A09714E29711BF4",
      X"731EFCACD21D053B0BDEFC521D514E7CAC8668724971E4934A22C971B0E63D50",
      X"30B3B4B858A76BDFABDF5510195B5EFC0668263C0696E9704DD14E28D9F11A08",
      -- Address 1024 to 1535
      X"BE03CADC52488CD3E0324873B44697EB20980C87C1304D7BF413E0CC873FFF01",
      X"19F1E4C73F55BB0B8A89256F2B7413B4B9F04D853B5FAB8B20676B2164931E57",
      X"EBDE5740CC869715EFD447C06668D95BA0334A23619B5E02C9246D7BA1CE7D50",
      X"5511B1B1B018F21CF80C78A696E8D8A73FAADCAD2F2A7643616439A46C873E57",
      X"D90FD54438595BF4463D511BA1311AF6BC52B7EB7545911B5FFE56BDFBF5EF7F",
      X"6697BEFD0590190F2B8B74121C531EA9714F819BF51018F3B412E29C52E236E8",
      X"E63CF859A53B0A7616BCF9A53AA29CF8580DD1E492E2C827954492E360CD7BA0",
      X"60666971B14ED7BE57BFAB2032B6BCF80DD04C780C2CD3E19AA29D50B2E33510",
      X"7C0794B9A59018A7C16590E6688D2ED74130190E83619AF6E827C0990F7FFE03",
      X"32E2C98F7FAA761714134BDE56E8266873E19B0A77BE561741CED642C8263DAE",
      X"D6BDAF80980D2F2BDEA98F80CDD0B2B740679446C236BD049249DAF6429DFBA0",
      X"AA2262636131E439F019F04C2DD1B14F7F54B95B5F54EC86C2C87248D90E7DAE",
      X"B31FAA8970B2B6E88D7AA236426334EC79A56ED7EB8A2237BEFCAD7AF7EBDFFF",
      X"CD2E7DFB0B20331E5616E92438A63C52E39E0237EB2130E66925C439A5C46DD0",
      X"CC79F0B34A7714EC2C78F34B754439F1B11AA2C925C5914F2A8924C7C19AF740",
      X"C0CCD2E2629DAE7DAF7E5741646C79F11BA099F01858A6C335453BA164C76B20",
      -- Address 1536 to 2047
      X"F90E28734B21314E83CB20CDD11A5DAE8360321C06C334EDD14F80331FFEFC07",
      X"65C4931FFF54ED2E282696BCADD04DD0E6C23715EE7CAD2E829CAD85904D7A5C",
      X"AD7B5F01311B5E56BC531F019BA1656F81CE288D846D7A092493B4ED853AF741",
      X"5545C4C6C262C873E033E0995AA2639FFEA872B7BEA8D80D8591E590B21DFA5C",
      X"673F5413E1646DD11BF5446D84C668D8F34ADDAED715456E7CF95BF5EED7BFFF",
      X"9A5DFAF61740663CAC2CD249704C79A4C63D056ED64360CCD34A88734A89DBA0",
      X"98F3E06795EE28D859F0E697EA8872E2633544934B8A239F5412498E8335EF81",
      X"8099A5C5C53A5DFB5EFDAE82C8D8F2E2374033E131B04C876B8A7642C98ED740",
      X"F21D50E69642629C0697419AA335BA5C07C164380C8669DAA39F00673EFCF90F",
      X"CA88273FFEA9DA5D504C2C795BA19BA0CD856F2ADCF95A5D04395B0B219BF4B8",
      X"5AF7BE026236BCAC78A73E023643CBDE029D511A09DBF412482669DB0B75EE83",
      X"AB8A888D85C590E7C067C033B544C73EFD51E56E7D51B11B0A23CB21653BF4B9",
      X"CF7EA826C2C9DAA237EA89DA088DD1B0E795BA5DAF2B8ADCF8F2B7EADDAF7FFF",
      X"35BBF4ED2F80CC785859A493E098F2488D7B0ADCAC87C098A79510E79412B741",
      X"30E7C1CF2ADD51B0B3E0CD2FD511E5C4C76A88269714473EA924921C076BDE03",
      X"00334B8B8B75BAF6BDFA5D0591B1E5C56F8066C26360990ED714ED84921DAF81"
);

--------------------------------------------------------
--      IMPLEMENTATION
--------------------------------------------------------
begin
-- Port A read
process(CLKA, ADDRA)
variable ROWA: integer range 0 to (2**(ADDR_WIDTH-5))-1 := 0;
variable COLA: integer range 0 to 255 := 0;
variable ADDRAL: std_logic_vector(7 downto 0) := (others => '0');
begin
	ROWA := to_integer(unsigned(not ADDRA(ADDRA'left downto 5)));	-- 32 bytes per row, reading from top to bottom
	ADDRAL := ADDRA(4 downto 0) & "000";	-- selected byte in a row, reading from right to left
	COLA := to_integer(unsigned(ADDRAL));	

	if rising_edge(CLKA) then
		if(CSA = '1') then
			DOA_local <= ROM(ROWA)(COLA+7 downto COLA);
		else
			DOA_local <= (others => '0');
		end if;
	end if;
end process;

-- tri-state output
DOA <= DOA_local when (CSA = '1') and (OEA = '1') else (others => 'Z');
 

-- Port B read
process(CLKB, ADDRB)
variable ROWB: integer range 0 to (2**(ADDR_WIDTH-5))-1 := 0;
variable COLB: integer range 0 to 255 := 0;
variable ADDRBL: std_logic_vector(7 downto 0) := (others => '0');
begin
	ROWB := to_integer(unsigned(not ADDRB(ADDRB'left downto 5)));	-- 32 bytes per row, reading from top to bottom
	ADDRBL := ADDRB(4 downto 0) & "000";
	COLB := to_integer(unsigned(ADDRBL));	


	if rising_edge(CLKB) then
		if(CSB = '1') then
			DOB_local <= ROM(ROWB)(COLB+7 downto COLB);
		else
			DOB_local <= (others => '0');
		end if;
	end if;
end process;

-- tri-state output
DOB <= DOB_local when (CSB = '1') and (OEB = '1') else (others => 'Z');

end Behavioral;
