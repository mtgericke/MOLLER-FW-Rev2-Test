-------------------------------------------------------------
-- Filename:  CRC32_LUT1cd.VHD
-- Authors: 
-- 	from http://www.xilinx.com/support/documentation/sw_manuals/xilinx14_4/xst_v6s6.pdf  p262
--		Alain Zarembowitch / MSS
-- Version: Rev 0
-- Last modified: 12/13/17
-- Inheritance: 	ROM1.vhd 8/24/16
--
-- description:  synthesizable generic dual port ROM containing two tables of 256 CRC32s values each
-- (called LUT1c and LUT1d)
-- The tables are generated by the Java application crc32tables in the /java folder
-- LUT1c computes the CRC32s for inputs in the form 00 x 00 00
-- LUT1d computes the CRC32s for inputs in the form y 00 00 00, where y is the MSB
-- Data bit order: MSb of MSB is first sent/received
-- Note: the returned crc values are NOT inverted and NOT reflected left-right. They are as they would appear
-- when generated by a standard LFSR
---------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity CRC32_LUT1cd is
	 Generic (
		DATA_WIDTH: integer := 32;	
		ADDR_WIDTH: integer := 9
	);
    Port ( 
	    -- Port A
		ADDRA  : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
			-- LUT1c at addresses 0 - 255
			-- LUT1d at addresses 256 - 511
		DOA  : out std_logic_vector(DATA_WIDTH-1 downto 0);

		-- Port B
		ADDRB  : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
			-- LUT1c at addresses 0 - 255
			-- LUT1d at addresses 256 - 511
		DOB  : out std_logic_vector(DATA_WIDTH-1 downto 0)
		);
end entity;

architecture Behavioral of CRC32_LUT1cd is
--------------------------------------------------------
--     SIGNALS
--------------------------------------------------------
-- inferred rom
signal DOA_local: std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
signal DOB_local: std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
type ROM_TYPE is array ( (2**ADDR_WIDTH)-1 downto 0 ) of std_logic_vector(DATA_WIDTH-1 downto 0);
-- IMPORTANT ORDER INFORMATION: the table below is read from bottom to top and right to left. Thus
-- to restore a common-sense order, address bits are inverted.
constant ROM : ROM_TYPE := (
-- LUT1c
x"00000000", x"01D8AC87", x"03B1590E", x"0269F589", x"0762B21C", x"06BA1E9B", x"04D3EB12", x"050B4795", 
x"0EC56438", x"0F1DC8BF", x"0D743D36", x"0CAC91B1", x"09A7D624", x"087F7AA3", x"0A168F2A", x"0BCE23AD", 
x"1D8AC870", x"1C5264F7", x"1E3B917E", x"1FE33DF9", x"1AE87A6C", x"1B30D6EB", x"19592362", x"18818FE5", 
x"134FAC48", x"129700CF", x"10FEF546", x"112659C1", x"142D1E54", x"15F5B2D3", x"179C475A", x"1644EBDD", 
x"3B1590E0", x"3ACD3C67", x"38A4C9EE", x"397C6569", x"3C7722FC", x"3DAF8E7B", x"3FC67BF2", x"3E1ED775", 
x"35D0F4D8", x"3408585F", x"3661ADD6", x"37B90151", x"32B246C4", x"336AEA43", x"31031FCA", x"30DBB34D", 
x"269F5890", x"2747F417", x"252E019E", x"24F6AD19", x"21FDEA8C", x"2025460B", x"224CB382", x"23941F05", 
x"285A3CA8", x"2982902F", x"2BEB65A6", x"2A33C921", x"2F388EB4", x"2EE02233", x"2C89D7BA", x"2D517B3D", 
x"762B21C0", x"77F38D47", x"759A78CE", x"7442D449", x"714993DC", x"70913F5B", x"72F8CAD2", x"73206655", 
x"78EE45F8", x"7936E97F", x"7B5F1CF6", x"7A87B071", x"7F8CF7E4", x"7E545B63", x"7C3DAEEA", x"7DE5026D", 
x"6BA1E9B0", x"6A794537", x"6810B0BE", x"69C81C39", x"6CC35BAC", x"6D1BF72B", x"6F7202A2", x"6EAAAE25", 
x"65648D88", x"64BC210F", x"66D5D486", x"670D7801", x"62063F94", x"63DE9313", x"61B7669A", x"606FCA1D", 
x"4D3EB120", x"4CE61DA7", x"4E8FE82E", x"4F5744A9", x"4A5C033C", x"4B84AFBB", x"49ED5A32", x"4835F6B5", 
x"43FBD518", x"4223799F", x"404A8C16", x"41922091", x"44996704", x"4541CB83", x"47283E0A", x"46F0928D", 
x"50B47950", x"516CD5D7", x"5305205E", x"52DD8CD9", x"57D6CB4C", x"560E67CB", x"54679242", x"55BF3EC5", 
x"5E711D68", x"5FA9B1EF", x"5DC04466", x"5C18E8E1", x"5913AF74", x"58CB03F3", x"5AA2F67A", x"5B7A5AFD", 
x"EC564380", x"ED8EEF07", x"EFE71A8E", x"EE3FB609", x"EB34F19C", x"EAEC5D1B", x"E885A892", x"E95D0415", 
x"E29327B8", x"E34B8B3F", x"E1227EB6", x"E0FAD231", x"E5F195A4", x"E4293923", x"E640CCAA", x"E798602D", 
x"F1DC8BF0", x"F0042777", x"F26DD2FE", x"F3B57E79", x"F6BE39EC", x"F766956B", x"F50F60E2", x"F4D7CC65", 
x"FF19EFC8", x"FEC1434F", x"FCA8B6C6", x"FD701A41", x"F87B5DD4", x"F9A3F153", x"FBCA04DA", x"FA12A85D", 
x"D743D360", x"D69B7FE7", x"D4F28A6E", x"D52A26E9", x"D021617C", x"D1F9CDFB", x"D3903872", x"D24894F5", 
x"D986B758", x"D85E1BDF", x"DA37EE56", x"DBEF42D1", x"DEE40544", x"DF3CA9C3", x"DD555C4A", x"DC8DF0CD", 
x"CAC91B10", x"CB11B797", x"C978421E", x"C8A0EE99", x"CDABA90C", x"CC73058B", x"CE1AF002", x"CFC25C85", 
x"C40C7F28", x"C5D4D3AF", x"C7BD2626", x"C6658AA1", x"C36ECD34", x"C2B661B3", x"C0DF943A", x"C10738BD", 
x"9A7D6240", x"9BA5CEC7", x"99CC3B4E", x"981497C9", x"9D1FD05C", x"9CC77CDB", x"9EAE8952", x"9F7625D5", 
x"94B80678", x"9560AAFF", x"97095F76", x"96D1F3F1", x"93DAB464", x"920218E3", x"906BED6A", x"91B341ED", 
x"87F7AA30", x"862F06B7", x"8446F33E", x"859E5FB9", x"8095182C", x"814DB4AB", x"83244122", x"82FCEDA5", 
x"8932CE08", x"88EA628F", x"8A839706", x"8B5B3B81", x"8E507C14", x"8F88D093", x"8DE1251A", x"8C39899D", 
x"A168F2A0", x"A0B05E27", x"A2D9ABAE", x"A3010729", x"A60A40BC", x"A7D2EC3B", x"A5BB19B2", x"A463B535", 
x"AFAD9698", x"AE753A1F", x"AC1CCF96", x"ADC46311", x"A8CF2484", x"A9178803", x"AB7E7D8A", x"AAA6D10D", 
x"BCE23AD0", x"BD3A9657", x"BF5363DE", x"BE8BCF59", x"BB8088CC", x"BA58244B", x"B831D1C2", x"B9E97D45", 
x"B2275EE8", x"B3FFF26F", x"B19607E6", x"B04EAB61", x"B545ECF4", x"B49D4073", x"B6F4B5FA", x"B72C197D", 
-- LUT1d
x"00000000", x"DC6D9AB7", x"BC1A28D9", x"6077B26E", x"7CF54C05", x"A098D6B2", x"C0EF64DC", x"1C82FE6B", 
x"F9EA980A", x"258702BD", x"45F0B0D3", x"999D2A64", x"851FD40F", x"59724EB8", x"3905FCD6", x"E5686661", 
x"F7142DA3", x"2B79B714", x"4B0E057A", x"97639FCD", x"8BE161A6", x"578CFB11", x"37FB497F", x"EB96D3C8", 
x"0EFEB5A9", x"D2932F1E", x"B2E49D70", x"6E8907C7", x"720BF9AC", x"AE66631B", x"CE11D175", x"127C4BC2", 
x"EAE946F1", x"3684DC46", x"56F36E28", x"8A9EF49F", x"961C0AF4", x"4A719043", x"2A06222D", x"F66BB89A", 
x"1303DEFB", x"CF6E444C", x"AF19F622", x"73746C95", x"6FF692FE", x"B39B0849", x"D3ECBA27", x"0F812090", 
x"1DFD6B52", x"C190F1E5", x"A1E7438B", x"7D8AD93C", x"61082757", x"BD65BDE0", x"DD120F8E", x"017F9539", 
x"E417F358", x"387A69EF", x"580DDB81", x"84604136", x"98E2BF5D", x"448F25EA", x"24F89784", x"F8950D33", 
x"D1139055", x"0D7E0AE2", x"6D09B88C", x"B164223B", x"ADE6DC50", x"718B46E7", x"11FCF489", x"CD916E3E", 
x"28F9085F", x"F49492E8", x"94E32086", x"488EBA31", x"540C445A", x"8861DEED", x"E8166C83", x"347BF634", 
x"2607BDF6", x"FA6A2741", x"9A1D952F", x"46700F98", x"5AF2F1F3", x"869F6B44", x"E6E8D92A", x"3A85439D", 
x"DFED25FC", x"0380BF4B", x"63F70D25", x"BF9A9792", x"A31869F9", x"7F75F34E", x"1F024120", x"C36FDB97", 
x"3BFAD6A4", x"E7974C13", x"87E0FE7D", x"5B8D64CA", x"470F9AA1", x"9B620016", x"FB15B278", x"277828CF", 
x"C2104EAE", x"1E7DD419", x"7E0A6677", x"A267FCC0", x"BEE502AB", x"6288981C", x"02FF2A72", x"DE92B0C5", 
x"CCEEFB07", x"108361B0", x"70F4D3DE", x"AC994969", x"B01BB702", x"6C762DB5", x"0C019FDB", x"D06C056C", 
x"3504630D", x"E969F9BA", x"891E4BD4", x"5573D163", x"49F12F08", x"959CB5BF", x"F5EB07D1", x"29869D66", 
x"A6E63D1D", x"7A8BA7AA", x"1AFC15C4", x"C6918F73", x"DA137118", x"067EEBAF", x"660959C1", x"BA64C376", 
x"5F0CA517", x"83613FA0", x"E3168DCE", x"3F7B1779", x"23F9E912", x"FF9473A5", x"9FE3C1CB", x"438E5B7C", 
x"51F210BE", x"8D9F8A09", x"EDE83867", x"3185A2D0", x"2D075CBB", x"F16AC60C", x"911D7462", x"4D70EED5", 
x"A81888B4", x"74751203", x"1402A06D", x"C86F3ADA", x"D4EDC4B1", x"08805E06", x"68F7EC68", x"B49A76DF", 
x"4C0F7BEC", x"9062E15B", x"F0155335", x"2C78C982", x"30FA37E9", x"EC97AD5E", x"8CE01F30", x"508D8587", 
x"B5E5E3E6", x"69887951", x"09FFCB3F", x"D5925188", x"C910AFE3", x"157D3554", x"750A873A", x"A9671D8D", 
x"BB1B564F", x"6776CCF8", x"07017E96", x"DB6CE421", x"C7EE1A4A", x"1B8380FD", x"7BF43293", x"A799A824", 
x"42F1CE45", x"9E9C54F2", x"FEEBE69C", x"22867C2B", x"3E048240", x"E26918F7", x"821EAA99", x"5E73302E", 
x"77F5AD48", x"AB9837FF", x"CBEF8591", x"17821F26", x"0B00E14D", x"D76D7BFA", x"B71AC994", x"6B775323", 
x"8E1F3542", x"5272AFF5", x"32051D9B", x"EE68872C", x"F2EA7947", x"2E87E3F0", x"4EF0519E", x"929DCB29", 
x"80E180EB", x"5C8C1A5C", x"3CFBA832", x"E0963285", x"FC14CCEE", x"20795659", x"400EE437", x"9C637E80", 
x"790B18E1", x"A5668256", x"C5113038", x"197CAA8F", x"05FE54E4", x"D993CE53", x"B9E47C3D", x"6589E68A", 
x"9D1CEBB9", x"4171710E", x"2106C360", x"FD6B59D7", x"E1E9A7BC", x"3D843D0B", x"5DF38F65", x"819E15D2", 
x"64F673B3", x"B89BE904", x"D8EC5B6A", x"0481C1DD", x"18033FB6", x"C46EA501", x"A419176F", x"78748DD8", 
x"6A08C61A", x"B6655CAD", x"D612EEC3", x"0A7F7474", x"16FD8A1F", x"CA9010A8", x"AAE7A2C6", x"768A3871", 
x"93E25E10", x"4F8FC4A7", x"2FF876C9", x"F395EC7E", x"EF171215", x"337A88A2", x"530D3ACC", x"8F60A07B" 
	);

--------------------------------------------------------
--      IMPLEMENTATION
--------------------------------------------------------
begin

-- Port A read
DOA <= ROM(to_integer(unsigned(not ADDRA)));	-- see IMPORTANT ORDER INFORMATION above
 

-- Port B read
DOB <= ROM(to_integer(unsigned(not ADDRB)));	-- see IMPORTANT ORDER INFORMATION above

end Behavioral;
