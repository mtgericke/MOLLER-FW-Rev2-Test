-------------------------------------------------------------
-- Filename:  CRC32_LUT2cd.VHD
-- Authors: 
-- 	from http://www.xilinx.com/support/documentation/sw_manuals/xilinx14_4/xst_v6s6.pdf  p262
--		Alain Zarembowitch / MSS
-- Version: Rev 0
-- Last modified: 12/13/17
-- Inheritance: 	ROM1.vhd 8/24/16
--
-- description:  synthesizable generic dual port ROM containing two tables of 256 CRC32s values each
-- (called LUT2c and LUT2d)
-- The tables are generated by the Java application crc32tables in the /java folder
-- LUT1c computes the CRC32s for 64-BIT INPUT WORDS in the form 00 x 00 00 00 00 00 00 
-- LUT1d computes the CRC32s for 64-BIT INPUT WORDS in the form y 00 00 00 00 00 00 00, where y is the MSB
-- Data bit order: MSb of MSB is first sent/received
-- Note: the returned crc values are NOT inverted and NOT reflected left-right. They are as they would appear
-- when generated by a standard LFSR
---------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity CRC32_LUT2cd is
	 Generic (
		DATA_WIDTH: integer := 32;	
		ADDR_WIDTH: integer := 9
	);
    Port ( 
	    -- Port A
		ADDRA  : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
			-- LUT1c at addresses 0 - 255
			-- LUT1d at addresses 256 - 511
		DOA  : out std_logic_vector(DATA_WIDTH-1 downto 0);

		-- Port B
		ADDRB  : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
			-- LUT1c at addresses 0 - 255
			-- LUT1d at addresses 256 - 511
		DOB  : out std_logic_vector(DATA_WIDTH-1 downto 0)
		);
end entity;

architecture Behavioral of CRC32_LUT2cd is
--------------------------------------------------------
--     SIGNALS
--------------------------------------------------------
-- inferred rom
signal DOA_local: std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
signal DOB_local: std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
type ROM_TYPE is array ( (2**ADDR_WIDTH)-1 downto 0 ) of std_logic_vector(DATA_WIDTH-1 downto 0);
-- IMPORTANT ORDER INFORMATION: the table below is read from bottom to top and right to left. Thus
-- to restore a common-sense order, address bits are inverted.
constant ROM : ROM_TYPE := (
-- LUT2c
x"00000000", x"4F576811", x"9EAED022", x"D1F9B833", x"399CBDF3", x"76CBD5E2", x"A7326DD1", x"E86505C0", 
x"73397BE6", x"3C6E13F7", x"ED97ABC4", x"A2C0C3D5", x"4AA5C615", x"05F2AE04", x"D40B1637", x"9B5C7E26", 
x"E672F7CC", x"A9259FDD", x"78DC27EE", x"378B4FFF", x"DFEE4A3F", x"90B9222E", x"41409A1D", x"0E17F20C", 
x"954B8C2A", x"DA1CE43B", x"0BE55C08", x"44B23419", x"ACD731D9", x"E38059C8", x"3279E1FB", x"7D2E89EA", 
x"C824F22F", x"87739A3E", x"568A220D", x"19DD4A1C", x"F1B84FDC", x"BEEF27CD", x"6F169FFE", x"2041F7EF", 
x"BB1D89C9", x"F44AE1D8", x"25B359EB", x"6AE431FA", x"8281343A", x"CDD65C2B", x"1C2FE418", x"53788C09", 
x"2E5605E3", x"61016DF2", x"B0F8D5C1", x"FFAFBDD0", x"17CAB810", x"589DD001", x"89646832", x"C6330023", 
x"5D6F7E05", x"12381614", x"C3C1AE27", x"8C96C636", x"64F3C3F6", x"2BA4ABE7", x"FA5D13D4", x"B50A7BC5", 
x"9488F9E9", x"DBDF91F8", x"0A2629CB", x"457141DA", x"AD14441A", x"E2432C0B", x"33BA9438", x"7CEDFC29", 
x"E7B1820F", x"A8E6EA1E", x"791F522D", x"36483A3C", x"DE2D3FFC", x"917A57ED", x"4083EFDE", x"0FD487CF", 
x"72FA0E25", x"3DAD6634", x"EC54DE07", x"A303B616", x"4B66B3D6", x"0431DBC7", x"D5C863F4", x"9A9F0BE5", 
x"01C375C3", x"4E941DD2", x"9F6DA5E1", x"D03ACDF0", x"385FC830", x"7708A021", x"A6F11812", x"E9A67003", 
x"5CAC0BC6", x"13FB63D7", x"C202DBE4", x"8D55B3F5", x"6530B635", x"2A67DE24", x"FB9E6617", x"B4C90E06", 
x"2F957020", x"60C21831", x"B13BA002", x"FE6CC813", x"1609CDD3", x"595EA5C2", x"88A71DF1", x"C7F075E0", 
x"BADEFC0A", x"F589941B", x"24702C28", x"6B274439", x"834241F9", x"CC1529E8", x"1DEC91DB", x"52BBF9CA", 
x"C9E787EC", x"86B0EFFD", x"574957CE", x"181E3FDF", x"F07B3A1F", x"BF2C520E", x"6ED5EA3D", x"2182822C", 
x"2DD0EE65", x"62878674", x"B37E3E47", x"FC295656", x"144C5396", x"5B1B3B87", x"8AE283B4", x"C5B5EBA5", 
x"5EE99583", x"11BEFD92", x"C04745A1", x"8F102DB0", x"67752870", x"28224061", x"F9DBF852", x"B68C9043", 
x"CBA219A9", x"84F571B8", x"550CC98B", x"1A5BA19A", x"F23EA45A", x"BD69CC4B", x"6C907478", x"23C71C69", 
x"B89B624F", x"F7CC0A5E", x"2635B26D", x"6962DA7C", x"8107DFBC", x"CE50B7AD", x"1FA90F9E", x"50FE678F", 
x"E5F41C4A", x"AAA3745B", x"7B5ACC68", x"340DA479", x"DC68A1B9", x"933FC9A8", x"42C6719B", x"0D91198A", 
x"96CD67AC", x"D99A0FBD", x"0863B78E", x"4734DF9F", x"AF51DA5F", x"E006B24E", x"31FF0A7D", x"7EA8626C", 
x"0386EB86", x"4CD18397", x"9D283BA4", x"D27F53B5", x"3A1A5675", x"754D3E64", x"A4B48657", x"EBE3EE46", 
x"70BF9060", x"3FE8F871", x"EE114042", x"A1462853", x"49232D93", x"06744582", x"D78DFDB1", x"98DA95A0", 
x"B958178C", x"F60F7F9D", x"27F6C7AE", x"68A1AFBF", x"80C4AA7F", x"CF93C26E", x"1E6A7A5D", x"513D124C", 
x"CA616C6A", x"8536047B", x"54CFBC48", x"1B98D459", x"F3FDD199", x"BCAAB988", x"6D5301BB", x"220469AA", 
x"5F2AE040", x"107D8851", x"C1843062", x"8ED35873", x"66B65DB3", x"29E135A2", x"F8188D91", x"B74FE580", 
x"2C139BA6", x"6344F3B7", x"B2BD4B84", x"FDEA2395", x"158F2655", x"5AD84E44", x"8B21F677", x"C4769E66", 
x"717CE5A3", x"3E2B8DB2", x"EFD23581", x"A0855D90", x"48E05850", x"07B73041", x"D64E8872", x"9919E063", 
x"02459E45", x"4D12F654", x"9CEB4E67", x"D3BC2676", x"3BD923B6", x"748E4BA7", x"A577F394", x"EA209B85", 
x"970E126F", x"D8597A7E", x"09A0C24D", x"46F7AA5C", x"AE92AF9C", x"E1C5C78D", x"303C7FBE", x"7F6B17AF", 
x"E4376989", x"AB600198", x"7A99B9AB", x"35CED1BA", x"DDABD47A", x"92FCBC6B", x"43050458", x"0C526C49", 
-- LUT2d
x"00000000", x"5BA1DCCA", x"B743B994", x"ECE2655E", x"6A466E9F", x"31E7B255", x"DD05D70B", x"86A40BC1", 
x"D48CDD3E", x"8F2D01F4", x"63CF64AA", x"386EB860", x"BECAB3A1", x"E56B6F6B", x"09890A35", x"5228D6FF", 
x"ADD8A7CB", x"F6797B01", x"1A9B1E5F", x"413AC295", x"C79EC954", x"9C3F159E", x"70DD70C0", x"2B7CAC0A", 
x"79547AF5", x"22F5A63F", x"CE17C361", x"95B61FAB", x"1312146A", x"48B3C8A0", x"A451ADFE", x"FFF07134", 
x"5F705221", x"04D18EEB", x"E833EBB5", x"B392377F", x"35363CBE", x"6E97E074", x"8275852A", x"D9D459E0", 
x"8BFC8F1F", x"D05D53D5", x"3CBF368B", x"671EEA41", x"E1BAE180", x"BA1B3D4A", x"56F95814", x"0D5884DE", 
x"F2A8F5EA", x"A9092920", x"45EB4C7E", x"1E4A90B4", x"98EE9B75", x"C34F47BF", x"2FAD22E1", x"740CFE2B", 
x"262428D4", x"7D85F41E", x"91679140", x"CAC64D8A", x"4C62464B", x"17C39A81", x"FB21FFDF", x"A0802315", 
x"BEE0A442", x"E5417888", x"09A31DD6", x"5202C11C", x"D4A6CADD", x"8F071617", x"63E57349", x"3844AF83", 
x"6A6C797C", x"31CDA5B6", x"DD2FC0E8", x"868E1C22", x"002A17E3", x"5B8BCB29", x"B769AE77", x"ECC872BD", 
x"13380389", x"4899DF43", x"A47BBA1D", x"FFDA66D7", x"797E6D16", x"22DFB1DC", x"CE3DD482", x"959C0848", 
x"C7B4DEB7", x"9C15027D", x"70F76723", x"2B56BBE9", x"ADF2B028", x"F6536CE2", x"1AB109BC", x"4110D576", 
x"E190F663", x"BA312AA9", x"56D34FF7", x"0D72933D", x"8BD698FC", x"D0774436", x"3C952168", x"6734FDA2", 
x"351C2B5D", x"6EBDF797", x"825F92C9", x"D9FE4E03", x"5F5A45C2", x"04FB9908", x"E819FC56", x"B3B8209C", 
x"4C4851A8", x"17E98D62", x"FB0BE83C", x"A0AA34F6", x"260E3F37", x"7DAFE3FD", x"914D86A3", x"CAEC5A69", 
x"98C48C96", x"C365505C", x"2F873502", x"7426E9C8", x"F282E209", x"A9233EC3", x"45C15B9D", x"1E608757", 
x"79005533", x"22A189F9", x"CE43ECA7", x"95E2306D", x"13463BAC", x"48E7E766", x"A4058238", x"FFA45EF2", 
x"AD8C880D", x"F62D54C7", x"1ACF3199", x"416EED53", x"C7CAE692", x"9C6B3A58", x"70895F06", x"2B2883CC", 
x"D4D8F2F8", x"8F792E32", x"639B4B6C", x"383A97A6", x"BE9E9C67", x"E53F40AD", x"09DD25F3", x"527CF939", 
x"00542FC6", x"5BF5F30C", x"B7179652", x"ECB64A98", x"6A124159", x"31B39D93", x"DD51F8CD", x"86F02407", 
x"26700712", x"7DD1DBD8", x"9133BE86", x"CA92624C", x"4C36698D", x"1797B547", x"FB75D019", x"A0D40CD3", 
x"F2FCDA2C", x"A95D06E6", x"45BF63B8", x"1E1EBF72", x"98BAB4B3", x"C31B6879", x"2FF90D27", x"7458D1ED", 
x"8BA8A0D9", x"D0097C13", x"3CEB194D", x"674AC587", x"E1EECE46", x"BA4F128C", x"56AD77D2", x"0D0CAB18", 
x"5F247DE7", x"0485A12D", x"E867C473", x"B3C618B9", x"35621378", x"6EC3CFB2", x"8221AAEC", x"D9807626", 
x"C7E0F171", x"9C412DBB", x"70A348E5", x"2B02942F", x"ADA69FEE", x"F6074324", x"1AE5267A", x"4144FAB0", 
x"136C2C4F", x"48CDF085", x"A42F95DB", x"FF8E4911", x"792A42D0", x"228B9E1A", x"CE69FB44", x"95C8278E", 
x"6A3856BA", x"31998A70", x"DD7BEF2E", x"86DA33E4", x"007E3825", x"5BDFE4EF", x"B73D81B1", x"EC9C5D7B", 
x"BEB48B84", x"E515574E", x"09F73210", x"5256EEDA", x"D4F2E51B", x"8F5339D1", x"63B15C8F", x"38108045", 
x"9890A350", x"C3317F9A", x"2FD31AC4", x"7472C60E", x"F2D6CDCF", x"A9771105", x"4595745B", x"1E34A891", 
x"4C1C7E6E", x"17BDA2A4", x"FB5FC7FA", x"A0FE1B30", x"265A10F1", x"7DFBCC3B", x"9119A965", x"CAB875AF", 
x"3548049B", x"6EE9D851", x"820BBD0F", x"D9AA61C5", x"5F0E6A04", x"04AFB6CE", x"E84DD390", x"B3EC0F5A", 
x"E1C4D9A5", x"BA65056F", x"56876031", x"0D26BCFB", x"8B82B73A", x"D0236BF0", x"3CC10EAE", x"6760D264"
	);

--------------------------------------------------------
--      IMPLEMENTATION
--------------------------------------------------------
begin

-- Port A read
DOA <= ROM(to_integer(unsigned(not ADDRA)));	-- see IMPORTANT ORDER INFORMATION above
 

-- Port B read
DOB <= ROM(to_integer(unsigned(not ADDRB)));	-- see IMPORTANT ORDER INFORMATION above

end Behavioral;
