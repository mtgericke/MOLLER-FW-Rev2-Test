-------------------------------------------------------------
-- MSS copyright 2017-2020
-- Filename:  COM1800_TOP.VHD
-- Authors:
--		Alain Zarembowitch / MSS
-- Version: Rev 4
-- Last modified: 10/25/20
-- Inheritance: 	n/a
--
-- description:  Top level for COM-1800 FPGA development platform
-- Includes only 10G Ethernet MAC + XAUI wrapper (using Xilinx transceiver wizzard 3.6 IP core)
-- For other COM-1800 features, download the com-1800 vhdl code template from
-- https://comblock.com/download.html#Latest_FPGA_firmware
--
-- In the case of Xilinx Artix -1 speed grade (slowest), better timing may be obtain by setting
--Project Settings | Synthesis | Options | keep equivalent registers, no resource sharing
---------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
Library UNISIM;
use UNISIM.vcomponents.all;

entity COM1800_TOP is
	generic (
		OPTION: std_logic_vector(7 downto 0) := x"20";    -- '-'    -- N/A
		REVISION: std_logic_vector(7 downto 0) := x"34";    -- '4'
		--// FPGA option and revision (ASCII format '0' = x30, 'A' = x41)
		-- These two ASCII characters appear in the Comblock Control Center.
		-- Helpful in identifying which firmware version is currently running in the FPGA.
		-- Select internal vs external frequency reference option.
		-- REMINDER: do change the .xdc file according to the option selection -A or -B
		SIMULATION: std_logic := '0'
		-- 1 during simulation, 0 for release
	);
    Port (
		--GLOBAL CLOCKS
	   CLKREF_TCXO : in std_logic;
			-- 19.2MHz reference clock. Generated by the VCTCXO on this board.
		CLKREF_EXT: in std_logic;
			-- external (higher-stability) frequency reference via J9 SMA connector ("EXT REF")

		-- 4 XAUI pairs for connection to 10GBASE Ethernet PHY
		MGTREFCLK0N: in std_logic;	-- 156.25 MHz differential clock
		MGTREFCLK0P: in std_logic;	-- requires installation of U10 156.26 MHz SMT oscillator
		XAUI_TX_L0_P : out std_logic;	-- @ 3.125 Gbits/s
		XAUI_TX_L0_N : out std_logic;
		XAUI_TX_L1_P : out std_logic;
		XAUI_TX_L1_N : out std_logic;
		XAUI_TX_L2_P : out std_logic;
		XAUI_TX_L2_N : out std_logic;
		XAUI_TX_L3_P : out std_logic;
		XAUI_TX_L3_N : out std_logic;
		XAUI_RX_L0_P : in std_logic;
		XAUI_RX_L0_N : in std_logic;
		XAUI_RX_L1_P : in std_logic;
		XAUI_RX_L1_N : in std_logic;
		XAUI_RX_L2_P : in std_logic;
		XAUI_RX_L2_N : in std_logic;
		XAUI_RX_L3_P : in std_logic;
		XAUI_RX_L3_N : in std_logic;

		--// Left connector, 98 pin PCIe female connector.
		-- Pins B5,B20,B31,B42 reserved for Ground
		-- Pins A49/B49 reserved for ComBlock Monitoring and Control.
		-- Place B13 in high-impedance when using the 12-bit DAC or vice versa.
		-- Hardware connects LEFT_CONNECTOR_A(38:32) with LEFT_CONNECTOR_B2(16:10)
		LEFT_CONNECTOR_A: inout std_logic_vector(38 downto 1);
		LEFT_CONNECTOR_B1: inout std_logic_vector(4 downto 1);
		LEFT_CONNECTOR_B2: inout std_logic_vector(16 downto 6);

		--// Right connector: 98 pin PCIe female connector.
		-- Pins B5,B20,B31,B42 reserved for Ground
		-- Pins A49/B49 reserved for ComBlock Monitoring and Control.
		-- Connector pins A39 - A48, B40,B41,B43-B48 can be used by
		-- re-routing LEFT_CONNECTOR signals using a resistor array (requires soldering)
		-- See schematics for details.
		RIGHT_CONNECTOR_A: inout std_logic_vector(38 downto 1);
		RIGHT_CONNECTOR_B1: inout std_logic_vector(4 downto 1);
		RIGHT_CONNECTOR_B2: inout std_logic_vector(19 downto 6);
		RIGHT_CONNECTOR_B3: inout std_logic_vector(30 downto 21);
		RIGHT_CONNECTOR_B4: inout std_logic_vector(39 downto 32);



		--// Monitoring & Control: ARM Cortex M3 microcontroller interface
		-- asynchronous bus (shared with NAND flash)
		-- set address at the rising edge of UC_WEB_IN when UC_CSIB_IN = '0' and UC_ALE_IN = '1'
		-- write data the rising edge of UC_WEB_IN when UC_CSIB_IN = '0'
		-- read data when  UC_CSIB_IN = '0' and UC_REB_IN = '0'
		UC_CSIB_IN: in std_logic;  -- chip select. active low.
		UC_ALE_IN: in std_logic;  -- address latch enable. active high.
		UC_REB_IN: in std_logic;  -- read enable #
		UC_WEB_IN: in std_logic;	-- write enable #
		UC_AD: inout std_logic_vector(7 downto 0)  -- shared address/data bus


			  );
end entity;

architecture Behavioral of COM1800_TOP is
--------------------------------------------------------
--      COMPONENTS
--------------------------------------------------------
-- Comment in/out components/drivers as needed

	COMPONENT CLKGEN7_MMCM_ADJ
	GENERIC (
		CLKFBOUT_MULT_F: real;
		CLKOUT0_DIVIDE_F: real;
		CLKIN1_PERIOD: real
    );
    PORT(
		CLK_IN1 : IN std_logic;
		CLK_OUT1 : OUT std_logic;
		PHASE_SHIFT_VAL: in std_logic_vector(7 downto 0);
		PHASE_SHIFT_TRIGGER_TOGGLE: in std_logic;
		INPUT_CLK_STOPPED : OUT std_logic;
		LOCKED : OUT std_logic;
		TP: OUT std_logic_vector(10 downto 1)
        );
    END COMPONENT;

component xaui_wrapper
port
(
    SOFT_RESET_TX_IN                        : in   std_logic;
    SOFT_RESET_RX_IN                        : in   std_logic;
    DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
    Q0_CLK0_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q0_CLK0_GTREFCLK_PAD_P_IN               : in   std_logic;
    Q0_CLK1_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q0_CLK1_GTREFCLK_PAD_P_IN               : in   std_logic;

    GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_DATA_VALID_IN                       : in   std_logic;
    GT1_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_DATA_VALID_IN                       : in   std_logic;
    GT2_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_DATA_VALID_IN                       : in   std_logic;
    GT3_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_DATA_VALID_IN                       : in   std_logic;

    GT0_TXUSRCLK_OUT                        : out  std_logic;
    GT0_TXUSRCLK2_OUT                       : out  std_logic;
    GT0_RXUSRCLK_OUT                        : out  std_logic;
    GT0_RXUSRCLK2_OUT                       : out  std_logic;

    GT1_TXUSRCLK_OUT                        : out  std_logic;
    GT1_TXUSRCLK2_OUT                       : out  std_logic;
    GT1_RXUSRCLK_OUT                        : out  std_logic;
    GT1_RXUSRCLK2_OUT                       : out  std_logic;

    GT2_TXUSRCLK_OUT                        : out  std_logic;
    GT2_TXUSRCLK2_OUT                       : out  std_logic;
    GT2_RXUSRCLK_OUT                        : out  std_logic;
    GT2_RXUSRCLK2_OUT                       : out  std_logic;

    GT3_TXUSRCLK_OUT                        : out  std_logic;
    GT3_TXUSRCLK2_OUT                       : out  std_logic;
    GT3_RXUSRCLK_OUT                        : out  std_logic;
    GT3_RXUSRCLK2_OUT                       : out  std_logic;

    --_________________________________________________________________________
    --GT0  (X0Y0)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt0_drpen_in                            : in   std_logic;
    gt0_drprdy_out                          : out  std_logic;
    gt0_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_eyescanreset_in                     : in   std_logic;
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    gt0_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    gt0_rxclkcorcnt_out                     : out  std_logic_vector(1 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxcharisk_out                       : out  std_logic_vector(1 downto 0);
    gt0_rxdisperr_out                       : out  std_logic_vector(1 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gtprxn_in                           : in   std_logic;
    gt0_gtprxp_in                           : in   std_logic;
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
    gt0_rxchanbondseq_out                   : out  std_logic;
    gt0_rxchbonden_in                       : in   std_logic;
    gt0_rxchbondi_in                        : in   std_logic_vector(3 downto 0);
    gt0_rxchbondlevel_in                    : in   std_logic_vector(2 downto 0);
    gt0_rxchbondmaster_in                   : in   std_logic;
    gt0_rxchbondo_out                       : out  std_logic_vector(3 downto 0);
    gt0_rxchbondslave_in                    : in   std_logic;
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
    gt0_rxchanisaligned_out                 : out  std_logic;
    gt0_rxchanrealign_out                   : out  std_logic;
    ------------ Receive Ports - RX Decision Feedback Equalizer(DFE) -----------
    gt0_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt0_rxlpmhfhold_in                      : in   std_logic;
    gt0_rxlpmhfovrden_in                    : in   std_logic;
    gt0_rxlpmlfhold_in                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    gt0_rxlpmreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt0_rxpolarity_in                       : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt0_txdata_in                           : in   std_logic_vector(15 downto 0);
    ------------------ Transmit Ports - TX 8B/10B Encoder Ports ----------------
    gt0_txcharisk_in                        : in   std_logic_vector(1 downto 0);
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt0_gtptxn_out                          : out  std_logic;
    gt0_gtptxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt0_txpolarity_in                       : in   std_logic;

    --GT1  (X0Y1)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt1_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt1_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt1_drpen_in                            : in   std_logic;
    gt1_drprdy_out                          : out  std_logic;
    gt1_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_eyescanreset_in                     : in   std_logic;
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    gt1_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    gt1_rxclkcorcnt_out                     : out  std_logic_vector(1 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt1_rxcharisk_out                       : out  std_logic_vector(1 downto 0);
    gt1_rxdisperr_out                       : out  std_logic_vector(1 downto 0);
    gt1_rxnotintable_out                    : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gtprxn_in                           : in   std_logic;
    gt1_gtprxp_in                           : in   std_logic;
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
    gt1_rxchanbondseq_out                   : out  std_logic;
    gt1_rxchbonden_in                       : in   std_logic;
    gt1_rxchbondi_in                        : in   std_logic_vector(3 downto 0);
    gt1_rxchbondlevel_in                    : in   std_logic_vector(2 downto 0);
    gt1_rxchbondmaster_in                   : in   std_logic;
    gt1_rxchbondo_out                       : out  std_logic_vector(3 downto 0);
    gt1_rxchbondslave_in                    : in   std_logic;
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
    gt1_rxchanisaligned_out                 : out  std_logic;
    gt1_rxchanrealign_out                   : out  std_logic;
    ------------ Receive Ports - RX Decision Feedback Equalizer(DFE) -----------
    gt1_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt1_rxlpmhfhold_in                      : in   std_logic;
    gt1_rxlpmhfovrden_in                    : in   std_logic;
    gt1_rxlpmlfhold_in                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt1_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    gt1_rxlpmreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt1_rxpolarity_in                       : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    gt1_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt1_txdata_in                           : in   std_logic_vector(15 downto 0);
    ------------------ Transmit Ports - TX 8B/10B Encoder Ports ----------------
    gt1_txcharisk_in                        : in   std_logic_vector(1 downto 0);
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt1_gtptxn_out                          : out  std_logic;
    gt1_gtptxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt1_txoutclkfabric_out                  : out  std_logic;
    gt1_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt1_txpolarity_in                       : in   std_logic;

    --GT2  (X0Y2)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt2_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt2_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt2_drpen_in                            : in   std_logic;
    gt2_drprdy_out                          : out  std_logic;
    gt2_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_eyescanreset_in                     : in   std_logic;
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    gt2_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    gt2_rxclkcorcnt_out                     : out  std_logic_vector(1 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt2_rxcharisk_out                       : out  std_logic_vector(1 downto 0);
    gt2_rxdisperr_out                       : out  std_logic_vector(1 downto 0);
    gt2_rxnotintable_out                    : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gtprxn_in                           : in   std_logic;
    gt2_gtprxp_in                           : in   std_logic;
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
    gt2_rxchanbondseq_out                   : out  std_logic;
    gt2_rxchbonden_in                       : in   std_logic;
    gt2_rxchbondi_in                        : in   std_logic_vector(3 downto 0);
    gt2_rxchbondlevel_in                    : in   std_logic_vector(2 downto 0);
    gt2_rxchbondmaster_in                   : in   std_logic;
    gt2_rxchbondo_out                       : out  std_logic_vector(3 downto 0);
    gt2_rxchbondslave_in                    : in   std_logic;
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
    gt2_rxchanisaligned_out                 : out  std_logic;
    gt2_rxchanrealign_out                   : out  std_logic;
    ------------ Receive Ports - RX Decision Feedback Equalizer(DFE) -----------
    gt2_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt2_rxlpmhfhold_in                      : in   std_logic;
    gt2_rxlpmhfovrden_in                    : in   std_logic;
    gt2_rxlpmlfhold_in                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt2_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    gt2_rxlpmreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt2_rxpolarity_in                       : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    gt2_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt2_txdata_in                           : in   std_logic_vector(15 downto 0);
    ------------------ Transmit Ports - TX 8B/10B Encoder Ports ----------------
    gt2_txcharisk_in                        : in   std_logic_vector(1 downto 0);
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt2_gtptxn_out                          : out  std_logic;
    gt2_gtptxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt2_txoutclkfabric_out                  : out  std_logic;
    gt2_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt2_txpolarity_in                       : in   std_logic;

    --GT3  (X0Y3)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt3_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt3_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt3_drpen_in                            : in   std_logic;
    gt3_drprdy_out                          : out  std_logic;
    gt3_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_eyescanreset_in                     : in   std_logic;
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    gt3_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    gt3_rxclkcorcnt_out                     : out  std_logic_vector(1 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(15 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt3_rxcharisk_out                       : out  std_logic_vector(1 downto 0);
    gt3_rxdisperr_out                       : out  std_logic_vector(1 downto 0);
    gt3_rxnotintable_out                    : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gtprxn_in                           : in   std_logic;
    gt3_gtprxp_in                           : in   std_logic;
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
    gt3_rxchanbondseq_out                   : out  std_logic;
    gt3_rxchbonden_in                       : in   std_logic;
    gt3_rxchbondi_in                        : in   std_logic_vector(3 downto 0);
    gt3_rxchbondlevel_in                    : in   std_logic_vector(2 downto 0);
    gt3_rxchbondmaster_in                   : in   std_logic;
    gt3_rxchbondo_out                       : out  std_logic_vector(3 downto 0);
    gt3_rxchbondslave_in                    : in   std_logic;
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
    gt3_rxchanisaligned_out                 : out  std_logic;
    gt3_rxchanrealign_out                   : out  std_logic;
    ------------ Receive Ports - RX Decision Feedback Equalizer(DFE) -----------
    gt3_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt3_rxlpmhfhold_in                      : in   std_logic;
    gt3_rxlpmhfovrden_in                    : in   std_logic;
    gt3_rxlpmlfhold_in                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt3_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    gt3_rxlpmreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt3_rxpolarity_in                       : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    gt3_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt3_txdata_in                           : in   std_logic_vector(15 downto 0);
    ------------------ Transmit Ports - TX 8B/10B Encoder Ports ----------------
    gt3_txcharisk_in                        : in   std_logic_vector(1 downto 0);
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt3_gtptxn_out                          : out  std_logic;
    gt3_gtptxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt3_txoutclkfabric_out                  : out  std_logic;
    gt3_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt3_txpolarity_in                       : in   std_logic;

    --____________________________COMMON PORTS________________________________
   GT0_PLL0RESET_OUT  : out std_logic;
         GT0_PLL0OUTCLK_OUT  : out std_logic;
         GT0_PLL0OUTREFCLK_OUT  : out std_logic;
         GT0_PLL0LOCK_OUT  : out std_logic;
         GT0_PLL0REFCLKLOST_OUT  : out std_logic;
         GT0_PLL1OUTCLK_OUT  : out std_logic;
         GT0_PLL1OUTREFCLK_OUT  : out std_logic;

          sysclk_in                               : in   std_logic

);

end component;

	COMPONENT XAUI2XGMII
	PORT(
		SYNC_RESET : IN std_logic;
		CLK : IN std_logic;
		XAUI_RXD : IN std_logic_vector(31 downto 0);
		XAUI_RXCHARISK : IN std_logic_vector(3 downto 0);
		XAUI_RXDISPERR : IN std_logic_vector(3 downto 0);
		XAUI_RXNOTINTABLE : IN std_logic_vector(3 downto 0);
		XGMII_RXD : OUT std_logic_vector(31 downto 0);
		XGMII_RXC : OUT std_logic_vector(3 downto 0)
		);
	END COMPONENT;

	COMPONENT XGMII2XAUI
	GENERIC (
		NBYTES: integer
    );
	PORT(
		SYNC_RESET : IN std_logic;
		CLK : IN std_logic;
		XGMII_TXD: in std_logic_vector(8*NBYTES-1 downto 0);
		XGMII_TXC: in std_logic_vector(NBYTES-1 downto 0);
		XAUI_TXD: out std_logic_vector(8*NBYTES-1 downto 0);
		XAUI_TXCHARISK: out std_logic_vector(NBYTES-1 downto 0);
		TP : OUT std_logic_vector(10 downto 1)
		);
	END COMPONENT;

	COMPONENT COM5501
	GENERIC (
		EXT_PHY_MDIO_ADDR: std_logic_vector(4 downto 0);
		RX_MTU: integer;
		RX_BUFFER: std_logic;
		RX_BUFFER_ADDR_NBITS: integer;
		TX_MTU: integer;
		TX_BUFFER: std_logic;
		TX_BUFFER_ADDR_NBITS: integer;
		MAC_CONTROL_PAUSE_ENABLE: std_logic;
		SIMULATION: std_logic
    );
	PORT(
		CLK : IN std_logic;
		SYNC_RESET : IN std_logic;
		CLK156g : IN std_logic;
		MAC_TX_CONFIG : IN std_logic_vector(7 downto 0);
		MAC_RX_CONFIG : IN std_logic_vector(7 downto 0);
		MAC_ADDR : IN std_logic_vector(47 downto 0);
		MAC_TX_DATA : IN std_logic_vector(63 downto 0);
		MAC_TX_DATA_VALID : IN std_logic_vector(7 downto 0);
		MAC_TX_EOF : IN std_logic;
		MAC_RX_CTS : IN std_logic;
		XGMII_RXD : IN std_logic_vector(63 downto 0);
		XGMII_RXC : IN std_logic_vector(7 downto 0);
		MDIO_IN : IN std_logic;
		MDIO_DIR : out std_logic;
		MAC_TX_CTS : OUT std_logic;
		MAC_RX_DATA : OUT std_logic_vector(63 downto 0);
		MAC_RX_DATA_VALID : OUT std_logic_vector(7 downto 0);
		MAC_RX_SOF : OUT std_logic;
		MAC_RX_EOF : OUT std_logic;
		MAC_RX_FRAME_VALID: out std_logic;
		XGMII_TXD : OUT std_logic_vector(63 downto 0);
		XGMII_TXC : OUT std_logic_vector(7 downto 0);
		RESET_N : OUT std_logic;
		MDC : OUT std_logic;
		MDIO_OUT : OUT std_logic;
		PHY_CONFIG_CHANGE : IN std_logic;
		PHY_RESET: in std_logic;
		TEST_MODE: in std_logic_vector(1 downto 0);
		POWER_DOWN: in std_logic;
		PHY_STATUS: out std_logic_vector(7 downto 0);
		PHY_STATUS2: out std_logic_vector(7 downto 0);
		PHY_ID : OUT std_logic_vector(15 downto 0);
		N_TX_FRAMES : OUT std_logic_vector(15 downto 0);
		N_RX_FRAMES : OUT std_logic_vector(15 downto 0);
		N_RX_BAD_CRCS : OUT std_logic_vector(15 downto 0);
		N_RX_FRAMES_TOO_SHORT : OUT std_logic_vector(15 downto 0);
		N_RX_FRAMES_TOO_LONG : OUT std_logic_vector(15 downto 0);
		N_RX_WRONG_ADDR : OUT std_logic_vector(15 downto 0);
		N_RX_LENGTH_ERRORS : OUT std_logic_vector(15 downto 0);
		RX_IPG: out std_logic_vector(7 downto 0);
		DEBUG1 : OUT std_logic_vector(63 downto 0);
		DEBUG2 : OUT std_logic_vector(63 downto 0);
		DEBUG3 : OUT std_logic_vector(63 downto 0);
		TP : OUT std_logic_vector(10 downto 1)
		);
	END COMPONENT;

	COMPONENT TIMER_4US
	GENERIC (
		CLK_FREQUENCY: integer
	);
	PORT(
		SYNC_RESET : IN std_logic;
		CLK : IN std_logic;
		TICK_4US : OUT std_logic;
		TICK_100MS: out std_logic
		);
	END COMPONENT;

 	COMPONENT DNA_ID
	GENERIC (
		CLK_FREQUENCY: integer
	);
	PORT(
		CLK : IN std_logic;
		SYNC_RESET : IN std_logic;
		ID_OUT : OUT std_logic_vector(56 downto 0) := (others => '0');
		ID_VALID_OUT : OUT std_logic;
		ID_SAMPLE_CLK_OUT : OUT std_logic
		);
	END COMPONENT;


--------------------------------------------------------
--     SIGNALS
--------------------------------------------------------
-- Suffix _D indicates a one CLK delayed version of the net with the same name
-- Suffix _X indicates an extended precision version of the net with the same name
-- Suffix _N indicates an inverted version of the net with the same name


--// CLOCKS, RESETS
signal CLKREF_TCXOg: std_logic := '0';
signal CLK10: std_logic := '0';
signal CLK10g: std_logic := '0';
signal CLK10g0: std_logic := '0';
signal CLK10g1: std_logic := '0';
signal CLK10_LOCKED: std_logic := '0';
signal CLK10_INPUT_CLK_STOPPED: std_logic := '0';
constant CLK_FREQUENCY: integer := 156; -- processing clock frequency CLK156g in MHz, as time reference
signal TICK_100MS: std_logic := '0';
signal TICK_1S: std_logic := '0';
signal TICK_1S_SHIFT: std_logic_vector(6 downto 0) := (others => '0');
signal TICK_4US: std_logic := '0';
signal TICK_100MS_CNTR: unsigned(3 downto 0) := (others => '0');
signal RESET_COUNTER: unsigned(23 downto 0) := x"000000";	-- initialize for simulations
	-- spans 2^23/10MHz = 838ms
signal RESET_STATE: integer range 0 to 2 := 0;
signal ASYNC_RESET: std_logic := '1';
signal SYNC_RESET_CLK156: std_logic := '0';
signal READY_FLAG_CLK156: std_logic := '0';

--//-- 10G ETHERNET XAUI ---------------------------------
signal CLK156: std_logic := '0';
signal CLK156g: std_logic := '0';
signal CLK156_LOCK: std_logic := '0';
signal CLK156_LOCK_D: std_logic := '0';
signal GT_TXUSERRDY: std_logic := '0';
signal XGMII_TXD : std_logic_vector(63 downto 0) := (others => '0');
signal XGMII_TXC : std_logic_vector(7 downto 0) := (others => '0');
signal XGMII_RXD1 : std_logic_vector(63 downto 0) := (others => '0');
signal XGMII_RXC1 : std_logic_vector(7 downto 0) := (others => '0');
signal XGMII_RXD : std_logic_vector(63 downto 0) := (others => '0');
signal XGMII_RXC : std_logic_vector(7 downto 0) := (others => '0');
signal XAUI_DEBUG: std_logic_vector(5 downto 0) := (others => '0');
signal XAUI_CONFIG: std_logic_vector(6 downto 0) := (others => '0');
signal gt0_txdata_in: std_logic_vector(15 downto 0) := (others => '0');
signal gt1_txdata_in: std_logic_vector(15 downto 0) := (others => '0');
signal gt2_txdata_in: std_logic_vector(15 downto 0) := (others => '0');
signal gt3_txdata_in: std_logic_vector(15 downto 0) := (others => '0');
signal gt0_rxdata_out: std_logic_vector(15 downto 0) := (others => '0');
signal gt1_rxdata_out: std_logic_vector(15 downto 0) := (others => '0');
signal gt2_rxdata_out: std_logic_vector(15 downto 0) := (others => '0');
signal gt3_rxdata_out: std_logic_vector(15 downto 0) := (others => '0');
signal GT0_PLL0RESET_OUT: std_logic := '0';
signal gt0_rxchbondo_out: std_logic_vector(3 downto 0) := (others => '0');
signal gt0_rxchanisaligned_out: std_logic := '0';
signal gt1_rxchanisaligned_out: std_logic := '0';
signal gt2_rxchanisaligned_out: std_logic := '0';
signal gt3_rxchanisaligned_out: std_logic := '0';
signal gt0_rxchanbondseq_out: std_logic := '0';
signal gt1_rxchanbondseq_out: std_logic := '0';
signal gt2_rxchanbondseq_out: std_logic := '0';
signal gt3_rxchanbondseq_out: std_logic := '0';
signal gt0_rxdisperr_out: std_logic_vector(1 downto 0) := (others => '0');
signal gt1_rxdisperr_out: std_logic_vector(1 downto 0) := (others => '0');
signal gt2_rxdisperr_out: std_logic_vector(1 downto 0) := (others => '0');
signal gt3_rxdisperr_out: std_logic_vector(1 downto 0) := (others => '0');
signal gt_rxpolarity_in: std_logic := '0';
signal gt_txpolarity_in: std_logic := '0';
signal gt0_rxcharisk_out: std_logic_vector(1 downto 0) := (others => '0');
signal gt1_rxcharisk_out: std_logic_vector(1 downto 0) := (others => '0');
signal gt2_rxcharisk_out: std_logic_vector(1 downto 0) := (others => '0');
signal gt3_rxcharisk_out: std_logic_vector(1 downto 0) := (others => '0');
signal gt0_rxnotintable_out: std_logic_vector(1 downto 0) := (others => '0');
signal gt1_rxnotintable_out: std_logic_vector(1 downto 0) := (others => '0');
signal gt2_rxnotintable_out: std_logic_vector(1 downto 0) := (others => '0');
signal gt3_rxnotintable_out: std_logic_vector(1 downto 0) := (others => '0');
signal gt0_txcharisk_in: std_logic_vector(1 downto 0) := (others => '0');
signal gt1_txcharisk_in: std_logic_vector(1 downto 0) := (others => '0');
signal gt2_txcharisk_in: std_logic_vector(1 downto 0) := (others => '0');
signal gt3_txcharisk_in: std_logic_vector(1 downto 0) := (others => '0');

--//-- XGMII INTERFACE ---------------------------------
signal XAUI_RXD: std_logic_vector(63 downto 0):= (others => '0');
signal XAUI_RXCHARISK: std_logic_vector(7 downto 0):= (others => '0');
signal XAUI_RXDISPERR: std_logic_vector(7 downto 0):= (others => '0');
signal XAUI_RXNOTINTABLE: std_logic_vector(7 downto 0):= (others => '0');
signal XAUI_TXD: std_logic_vector(63 downto 0):= (others => '0');
signal XAUI_TXCHARISK: std_logic_vector(7 downto 0):= (others => '0');
signal XAUI_TP: std_logic_vector(10 downto 1):= (others => '0');

--//-- ETHERNET MAC#1-----------------------------------
signal LAN1_MAC_ADDR: std_logic_vector(47 downto 0) := (others => '0');
signal LAN1_MDIO_IN: std_logic := '0';
signal LAN1_MDC: std_logic := '0';
signal LAN1_MDIO_OUT: std_logic := '0';
signal LAN1_MDIO_DIR: std_logic := '0';
signal LAN1_PHY_RESET: std_logic := '0';
signal LAN1_TEST_MODE: std_logic_vector(1 downto 0) := (others => '0');
signal LAN1_POWER_DOWN: std_logic := '0';
signal LAN1_PHY_ID: std_logic_vector(15 downto 0) := (others => '0');
signal LAN1_PHY_STATUS: std_logic_vector(7 downto 0) := (others => '0');
signal LAN1_PHY_STATUS2: std_logic_vector(7 downto 0) := (others => '0');
signal LAN1_N_RX_FRAMES: std_logic_vector(15 downto 0) := (others => '0');
signal LAN1_N_TX_FRAMES: std_logic_vector(15 downto 0) := (others => '0');
signal LAN1_MAC_TX_DATA: std_logic_vector(63 downto 0) := (others => '0');
signal LAN1_MAC_TX_DATA_VALID: std_logic_vector(7 downto 0) := (others => '0');
signal LAN1_MAC_TX_EOF: std_logic:= '0';
signal LAN1_MAC_TX_CTS: std_logic:= '0';
signal PHY_CONFIG_CHANGE: std_logic := '0';

signal DEBUG1: std_logic_vector(63 downto 0) := (others => '0');
signal DEBUG2: std_logic_vector(63 downto 0) := (others => '0');
signal DEBUG3: std_logic_vector(63 downto 0) := (others => '0');
signal LAN1_TP: std_logic_vector(10 downto 1) := (others => '0');
signal LAN1_N_RX_BAD_CRCS:  std_logic_vector(15 downto 0);
signal LAN1_RX_IPG: std_logic_vector(7 downto 0);

--// LAN/TCP-IP Interface for M&C (port 1028)
signal RX_LAN: std_logic_vector(7 downto 0) := (others => '0');
signal RX_LAN_SAMPLE_CLK_REQ: std_logic;
signal RX_LAN_BUFFER_EMPTY: std_logic := '1';
signal RX_LAN_BUFFER_EMPTY_D: std_logic := '1';
signal RX_LAN_BUFFER_EMPTY_D2: std_logic := '1';

--// Interface for M&C
signal SREG254_READ_TOGGLE_D: std_logic := '0';
signal SREG254_READ_TOGGLE_D2: std_logic := '0';

--//-- DNA Port ------------------------------------
signal DNA_ID_DATA: std_logic_vector(56 downto 0) := (others => '0');
signal DNA_ID_SAMPLE_CLK: std_logic := '0';

--// ARM co-processor interface
signal UC_WEBG: std_logic := '0';  -- WE# through global buffer
signal UC_REBG: std_logic := '0';	-- RE# through global buffer
signal UC_ADDRESS: unsigned(7 downto 0) := (others => '0');
signal UC_AD_LOCAL: std_logic_vector(7 downto 0) := (others => '0');
signal UC_RDN_D: std_logic := '0';
signal UC_RDN_D2: std_logic := '0';
signal CONFIG_CHANGE_TOGGLE: std_logic := '0';
signal CONFIG_CHANGE_TOGGLE_D: std_logic := '0';
signal CONFIG_CHANGE_TOGGLE_D2: std_logic := '0';
signal CONFIG_CHANGE_PULSE: std_logic := '0';

--// Control Registers
constant NCREGS: integer := 10;	-- number of control registers.
constant NCREG_IMIN: integer := 0;	-- starting at this index
constant NCREG_IMAX: integer := (NCREG_IMIN+NCREGS-1);
type SLV8xNCREGStype is array (integer range NCREG_IMIN to NCREG_IMAX) of std_logic_vector(7 downto 0);
signal CREG: SLV8xNCREGStype := (others => (others => '0'));
signal REG255: std_logic_vector(7 downto 0) := (others => '0');

--// User-defined status Registers (add as needed)
constant NSREGS: integer := 45;	-- number of status registers.
constant NSREG_IMIN: integer := 7;	-- starting at this index
constant NSREG_IMAX: integer := (NSREG_IMIN+NSREGS-1);
type SLV8xNSREGStype is array (integer range NSREG_IMIN to NSREG_IMAX) of std_logic_vector(7 downto 0);
signal SREG: SLV8xNSREGStype := (others => (others => '0'));
signal SREG7_READ_TOGGLE: std_logic := '0';
signal SREG7_READ_TOGGLE_D: std_logic := '0';
signal SREG7_READ_TOGGLE_D2: std_logic := '0';
signal LATCH_MONITORING_PULSE: std_logic := '0';
signal SREG254_READ_TOGGLE: std_logic := '0';


signal TEST_CLK_CNTR: unsigned(15 downto 0) := (others => '0');
--------------------------------------------------------
--      IMPLEMENTATION
--------------------------------------------------------
begin
--//--------------------------------------------------------------------------
--// CLOCKS, RESETS
--//--------------------------------------------------------------------------
-- Frequency plan:
-- 19.2 MHz TCXO or 10 MHz external -> 160 MHz (one of several possible CLK_TX)
-- -> 125 MHz with multiple phases (CLK_P, Ethernet LAN PHY)
-- 156.25 MHz processing clock from oscillator on the board.

SIM_001: if(SIMULATION = '1') generate
	 -- 10 MHz
    process
    begin
        CLK10g <= '0';
        wait for 50 ns;
        CLK10g <= '1';
        wait for 50 ns;
    end process;
	 CLK10_LOCKED <= '1';
	 CLK10_INPUT_CLK_STOPPED <= '0';

    -- 19.2 MHz
    process
    begin
        CLKREF_TCXOg <= '0';
        wait for 26.04 ns;
        CLKREF_TCXOg <= '1';
        wait for 26.04 ns;
    end process;

end generate;

REF_CLK_GEN_002: if(SIMULATION = '0') generate
   BUFG_001: BUFG port map(I => CLKREF_TCXO, O=> CLKREF_TCXOg);
   BUFG_002: BUFG port map (I => CLKREF_EXT, O => CLK10g1);

    -- generate alternative 10MHz clock from the always-present 19.2MHz TCXO clock
     CLKGEN7C_001: CLKGEN7_MMCM_ADJ
    GENERIC MAP(
		CLKFBOUT_MULT_F => 50.000,
		CLKOUT0_DIVIDE_F => 96.000,
		CLKIN1_PERIOD => 52.083
    )
    PORT MAP(
		CLK_IN1 => CLKREF_TCXOg,    -- 19.2 MHz TCXO clock
		CLK_OUT1 => CLK10g0,    -- 10 MHz global
		PHASE_SHIFT_VAL => x"00",
		PHASE_SHIFT_TRIGGER_TOGGLE => '0',
		INPUT_CLK_STOPPED => CLK10_INPUT_CLK_STOPPED,
		LOCKED => CLK10_LOCKED,
		TP => open
    );

	-- select reference clock
	BUFGMUX_001 : BUFGMUX
	port map (
		O => CLK10g,   -- 1-bit output: Clock output
		I0 => CLK10g0, -- 1-bit input: Clock input (S=0)
		I1 => CLK10g1, -- 1-bit input: Clock input (S=1)
		S => CREG(0)(7)    -- 1-bit input: Clock select
	);

end generate;

-- report clocks status
SREG(9)(2 downto 0) <=  CLK156_LOCK & CLK10_LOCKED & (not CLK10_INPUT_CLK_STOPPED);

 -- Generate miscellaneous global clocks and resets from the
 -- external reference 10 MHz clock
 RESET_STATE_MACHINE_001: process(CLK10g)
 begin
	  if rising_edge(CLK10g) then
			-- PLL need time to lock. The reset of the application is still in reset
			if(RESET_COUNTER(17) = '0') and (SIMULATION = '0') then
				 -- wait a bit before asserting the PLL lock
				 RESET_COUNTER <= RESET_COUNTER + 1;
			elsif(RESET_COUNTER(5) = '0') and (SIMULATION = '1') then
				 -- make it short during simulations
				 -- wait a bit before asserting the PLL lock
				 RESET_COUNTER <= RESET_COUNTER + 1;
			elsif(RESET_STATE = 0) and (CLK10_LOCKED = '1') then
				 -- wait until the 10 MHz PLL are locked to generate a reset
				 -- Beware of circular logic (i.e. do not use CLK156_LOCK which may depend on ASYNC_RESET)
				 RESET_STATE <= 1;
			elsif(RESET_STATE = 1) and (CLK156_LOCK = '1') then
				RESET_STATE <= 2;
			end if;

			if(RESET_STATE = 0) then
				 ASYNC_RESET <= '1';
			else
				 ASYNC_RESET <= '0';
			end if;
	  end if;
 end process;

-- generate a reset synchronous with CLK156g
SYNC_RESET_CLK156_GEN: process(CLK156g)
begin
	if rising_edge(CLK156g) then
		CLK156_LOCK_D <= CLK156_LOCK;
	end if;
end process;
READY_FLAG_CLK156 <= CLK156_LOCK and CLK10_LOCKED;
SYNC_RESET_CLK156 <= '1' when (CLK156_LOCK = '1') and (CLK156_LOCK_D = '0') else
							CONFIG_CHANGE_PULSE and CLK156_LOCK;


	-- external input clock
BUFG_006: BUFG  port map (I=> UC_WEB_IN, O=> UC_WEBG);
	-- ARM WE#
BUFG_007: BUFG  port map (I=> UC_REB_IN, O=> UC_REBG);
	-- ARM RE#

-- 1s tick
TICK1S_001: TIMER_4US
GENERIC MAP(
	CLK_FREQUENCY => CLK_FREQUENCY
)
PORT MAP(
	SYNC_RESET => SYNC_RESET_CLK156,
	CLK => CLK156g,
	TICK_4US => TICK_4US,
	TICK_100MS => TICK_100MS
);

-- modulo-10 counter. 1s tick
TICK1S_002: process(CLK156g)
begin
	if rising_edge(CLK156g) then
		if(SYNC_RESET_CLK156 = '1') then
			TICK_100MS_CNTR <= "0000";
			TICK_1S <= '0';
		elsif(TICK_100MS = '1') then
			if(TICK_100MS_CNTR = 0) then
				TICK_100MS_CNTR <= "1001";
				TICK_1S <= '1';
			else
				TICK_100MS_CNTR <= TICK_100MS_CNTR - 1;
				TICK_1S <= '0';
			end if;
		else
			TICK_1S <= '0';
		end if;
	end if;
end process;

--//-- 10G ETHERNET XAUI ---------------------------------
-- Using Xilinx 7-series transceivers wizard (3.6) IP core
-- See Xilinx UG-482 for GTP configuration
-- See Xilinx PG168 for 7 series transceiver wizard configuration

GT_TXUSERRDY <= READY_FLAG_CLK156 and CLK156_LOCK and CLK10_LOCKED;
	--  drive TXUSERRDY High after these conditions are met:
	-- 1. All clocks used by the application including TXUSRCLK/TXUSRCLK2 are shown as stable or
	-- locked when the PLL or MMCM is used.
	-- 2. The user interface is ready to transmit data to the GTP transceiver



-- configure the GTP transceiver as follows:
-- Comma value: K28.5
   xaui_wrapper_i : xaui_wrapper
port map
(
    SOFT_RESET_TX_IN => '0',
    SOFT_RESET_RX_IN => '0',
    DONT_RESET_ON_DATA_ERROR_IN => '0',
    Q0_CLK0_GTREFCLK_PAD_N_IN => MGTREFCLK0N,   -- 156.25 MHz external oscillator
    Q0_CLK0_GTREFCLK_PAD_P_IN => MGTREFCLK0P,
    Q0_CLK1_GTREFCLK_PAD_N_IN => '0',
    Q0_CLK1_GTREFCLK_PAD_P_IN => '0',

     GT0_TX_FSM_RESET_DONE_OUT => open,
     GT0_RX_FSM_RESET_DONE_OUT => open,
     GT0_DATA_VALID_IN => '1',
     GT1_TX_FSM_RESET_DONE_OUT => open,
     GT1_RX_FSM_RESET_DONE_OUT => open,
     GT1_DATA_VALID_IN => '1',
     GT2_TX_FSM_RESET_DONE_OUT => open,
     GT2_RX_FSM_RESET_DONE_OUT => open,
     GT2_DATA_VALID_IN => '1',
     GT3_TX_FSM_RESET_DONE_OUT => open,
     GT3_RX_FSM_RESET_DONE_OUT => open,
     GT3_DATA_VALID_IN => '1',

     GT0_TXUSRCLK_OUT => CLK156,
     GT0_TXUSRCLK2_OUT => open,
     GT0_RXUSRCLK_OUT => open,
     GT0_RXUSRCLK2_OUT => open,

     GT1_TXUSRCLK_OUT => open,
     GT1_TXUSRCLK2_OUT => open,
     GT1_RXUSRCLK_OUT => open,
     GT1_RXUSRCLK2_OUT => open,

     GT2_TXUSRCLK_OUT => open,
     GT2_TXUSRCLK2_OUT => open,
     GT2_RXUSRCLK_OUT => open,
     GT2_RXUSRCLK2_OUT => open,

     GT3_TXUSRCLK_OUT => open,
     GT3_TXUSRCLK2_OUT => open,
     GT3_RXUSRCLK_OUT => open,
     GT3_RXUSRCLK2_OUT => open,

    --_________________________________________________________________________
    --GT0  (X0Y0)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
        gt0_drpaddr_in                  =>      (others => '0'),
        gt0_drpdi_in                    =>      (others => '0'),
        gt0_drpdo_out                   =>      open,
        gt0_drpen_in                    =>      '0',
        gt0_drprdy_out                  =>      open,
        gt0_drpwe_in                    =>      '0',
    --------------------- RX Initialization and Reset Ports --------------------
        gt0_eyescanreset_in             =>      '0',
        gt0_rxuserrdy_in                =>      READY_FLAG_CLK156,
    -------------------------- RX Margin Analysis Ports ------------------------
        gt0_eyescandataerror_out        =>      open,
        gt0_eyescantrigger_in           =>      '0',
    ------------------- Receive Ports - Clock Correction Ports -----------------
        gt0_rxclkcorcnt_out             =>      open,
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt0_rxdata_out                  =>      gt0_rxdata_out,
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt0_rxcharisk_out               =>      gt0_rxcharisk_out,
        gt0_rxdisperr_out               =>      gt0_rxdisperr_out,
        gt0_rxnotintable_out            =>      gt0_rxnotintable_out,
    ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt0_gtprxn_in                   =>      XAUI_RX_L0_N,
        gt0_gtprxp_in                   =>      XAUI_RX_L0_P,
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
        gt0_rxchanbondseq_out           =>      gt0_rxchanbondseq_out,
        gt0_rxchbonden_in               =>      '1',
        gt0_rxchbondi_in                =>      "0000",
        gt0_rxchbondlevel_in            =>      "001",	-- 3 slaves direct connection
        gt0_rxchbondmaster_in           =>      '1',	-- 0 master, 1,2,3 slave
        gt0_rxchbondo_out               =>      gt0_rxchbondo_out,
        gt0_rxchbondslave_in            =>      '0',
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
        gt0_rxchanisaligned_out         =>      gt0_rxchanisaligned_out,	-- meaningless???? this is the master
        gt0_rxchanrealign_out           =>      open,
    ------------ Receive Ports - RX Decision Feedback Equalizer(DFE) -----------
        gt0_dmonitorout_out             =>      open,
    -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt0_rxlpmhfhold_in              =>      '0',
        gt0_rxlpmhfovrden_in            =>      '0',
        gt0_rxlpmlfhold_in              =>      '0',
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt0_rxoutclkfabric_out          =>      open,
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt0_gtrxreset_in                =>      SYNC_RESET_CLK156,
        gt0_rxlpmreset_in               =>      '0',
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt0_rxpolarity_in               =>      gt_rxpolarity_in,
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt0_rxresetdone_out             =>      open,
    --------------------- TX Initialization and Reset Ports --------------------
        gt0_gttxreset_in                =>      SYNC_RESET_CLK156,
        gt0_txuserrdy_in                =>      GT_TXUSERRDY,
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt0_txdata_in                   =>      gt0_txdata_in,
    ------------------ Transmit Ports - TX 8B/10B Encoder Ports ----------------
        gt0_txcharisk_in                =>      gt0_txcharisk_in,
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
        gt0_gtptxn_out                  =>      XAUI_TX_L0_N,
        gt0_gtptxp_out                  =>      XAUI_TX_L0_P,
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt0_txoutclkfabric_out          =>      open,
        gt0_txoutclkpcs_out             =>      open,
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt0_txresetdone_out             =>      open,
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt0_txpolarity_in               =>      gt_txpolarity_in,

    --GT1  (X0Y1)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
        gt1_drpaddr_in                  =>      (others => '0'),
        gt1_drpdi_in                    =>      (others => '0'),
        gt1_drpdo_out                   =>      open,
        gt1_drpen_in                    =>      '0',
        gt1_drprdy_out                  =>      open,
        gt1_drpwe_in                    =>      '0',
    --------------------- RX Initialization and Reset Ports --------------------
        gt1_eyescanreset_in             =>      '0',
        gt1_rxuserrdy_in                =>      READY_FLAG_CLK156,
    -------------------------- RX Margin Analysis Ports ------------------------
        gt1_eyescandataerror_out        =>      open,
        gt1_eyescantrigger_in           =>      '0',
    ------------------- Receive Ports - Clock Correction Ports -----------------
        gt1_rxclkcorcnt_out             =>      open,
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt1_rxdata_out                  =>      gt1_rxdata_out,
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt1_rxcharisk_out               =>      gt1_rxcharisk_out,
        gt1_rxdisperr_out               =>      gt1_rxdisperr_out,
        gt1_rxnotintable_out            =>      gt1_rxnotintable_out,
    ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt1_gtprxn_in                   =>      XAUI_RX_L1_N,
        gt1_gtprxp_in                   =>      XAUI_RX_L1_P,
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
        gt1_rxchanbondseq_out           =>      gt1_rxchanbondseq_out,
        gt1_rxchbonden_in               =>      '1',
        gt1_rxchbondi_in                =>      gt0_rxchbondo_out,
        gt1_rxchbondlevel_in            =>      "000",	-- no more daisy chaining
        gt1_rxchbondmaster_in           =>      '0',
        gt1_rxchbondo_out               =>      open,
        gt1_rxchbondslave_in            =>      '1',	-- 0 master, 1,2,3 slave
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
        gt1_rxchanisaligned_out         =>      gt1_rxchanisaligned_out,
        gt1_rxchanrealign_out           =>      open,
    ------------ Receive Ports - RX Decision Feedback Equalizer(DFE) -----------
        gt1_dmonitorout_out             =>      open,
    -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt1_rxlpmhfhold_in              =>      '0',
        gt1_rxlpmhfovrden_in            =>      '0',
        gt1_rxlpmlfhold_in              =>      '0',
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt1_rxoutclkfabric_out          =>      open,
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt1_gtrxreset_in                =>      SYNC_RESET_CLK156,
        gt1_rxlpmreset_in               =>      '0',
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt1_rxpolarity_in               =>      gt_rxpolarity_in,
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt1_rxresetdone_out             =>      open,
    --------------------- TX Initialization and Reset Ports --------------------
        gt1_gttxreset_in                =>      SYNC_RESET_CLK156,
        gt1_txuserrdy_in                =>      GT_TXUSERRDY,
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt1_txdata_in                   =>      gt1_txdata_in,
    ------------------ Transmit Ports - TX 8B/10B Encoder Ports ----------------
        gt1_txcharisk_in                =>      gt1_txcharisk_in,
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
        gt1_gtptxn_out                  =>      XAUI_TX_L1_N,
        gt1_gtptxp_out                  =>      XAUI_TX_L1_P,
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt1_txoutclkfabric_out          =>      open,
        gt1_txoutclkpcs_out             =>      open,
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt1_txresetdone_out             =>      open,
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt1_txpolarity_in               =>      gt_txpolarity_in,

    --GT2  (X0Y2)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
        gt2_drpaddr_in                  =>      (others => '0'),
        gt2_drpdi_in                    =>      (others => '0'),
        gt2_drpdo_out                   =>      open,
        gt2_drpen_in                    =>      '0',
        gt2_drprdy_out                  =>      open,
        gt2_drpwe_in                    =>      '0',
    --------------------- RX Initialization and Reset Ports --------------------
        gt2_eyescanreset_in             =>      '0',
        gt2_rxuserrdy_in                =>      READY_FLAG_CLK156,
    -------------------------- RX Margin Analysis Ports ------------------------
        gt2_eyescandataerror_out        =>      open,
        gt2_eyescantrigger_in           =>      '0',
    ------------------- Receive Ports - Clock Correction Ports -----------------
        gt2_rxclkcorcnt_out             =>      open,
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt2_rxdata_out                  =>     gt2_rxdata_out,
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt2_rxcharisk_out               =>      gt2_rxcharisk_out,
        gt2_rxdisperr_out               =>      gt2_rxdisperr_out,
        gt2_rxnotintable_out            =>      gt2_rxnotintable_out,
    ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt2_gtprxn_in                   =>      XAUI_RX_L2_N,
        gt2_gtprxp_in                   =>      XAUI_RX_L2_P,
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
        gt2_rxchanbondseq_out           =>      gt2_rxchanbondseq_out,
        gt2_rxchbonden_in               =>      '1',
        gt2_rxchbondi_in                =>      gt0_rxchbondo_out,
        gt2_rxchbondlevel_in            =>      "000",	-- no more daisy chaining
        gt2_rxchbondmaster_in           =>      '0',
        gt2_rxchbondo_out               =>      open,
        gt2_rxchbondslave_in            =>      '1',	-- 0 master, 1,2,3 slave
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
        gt2_rxchanisaligned_out         =>      gt2_rxchanisaligned_out,
        gt2_rxchanrealign_out           =>      open,
    ------------ Receive Ports - RX Decision Feedback Equalizer(DFE) -----------
        gt2_dmonitorout_out             =>      open,
    -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt2_rxlpmhfhold_in              =>      '0',
        gt2_rxlpmhfovrden_in            =>      '0',
        gt2_rxlpmlfhold_in              =>      '0',
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt2_rxoutclkfabric_out          =>      open,
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt2_gtrxreset_in                =>      SYNC_RESET_CLK156,
        gt2_rxlpmreset_in               =>      '0',
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt2_rxpolarity_in               =>      gt_rxpolarity_in,
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt2_rxresetdone_out             =>      open,
    --------------------- TX Initialization and Reset Ports --------------------
        gt2_gttxreset_in                =>      SYNC_RESET_CLK156,
        gt2_txuserrdy_in                =>      GT_TXUSERRDY,
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt2_txdata_in                   =>      gt2_txdata_in,
    ------------------ Transmit Ports - TX 8B/10B Encoder Ports ----------------
        gt2_txcharisk_in                =>      gt2_txcharisk_in,
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
        gt2_gtptxn_out                  =>      XAUI_TX_L2_N,
        gt2_gtptxp_out                  =>      XAUI_TX_L2_P,
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt2_txoutclkfabric_out          =>      open,
        gt2_txoutclkpcs_out             =>      open,
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt2_txresetdone_out             =>      open,
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt2_txpolarity_in               =>      gt_txpolarity_in,

    --GT3  (X0Y3)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
        gt3_drpaddr_in                  =>      (others => '0'),
        gt3_drpdi_in                    =>      (others => '0'),
        gt3_drpdo_out                   =>      open,
        gt3_drpen_in                    =>      '0',
        gt3_drprdy_out                  =>      open,
        gt3_drpwe_in                    =>      '0',
    --------------------- RX Initialization and Reset Ports --------------------
        gt3_eyescanreset_in             =>      '0',
        gt3_rxuserrdy_in                =>      READY_FLAG_CLK156,
    -------------------------- RX Margin Analysis Ports ------------------------
        gt3_eyescandataerror_out        =>      open,
        gt3_eyescantrigger_in           =>      '0',
    ------------------- Receive Ports - Clock Correction Ports -----------------
        gt3_rxclkcorcnt_out             =>      open,
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt3_rxdata_out                  =>      gt3_rxdata_out,
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt3_rxcharisk_out               =>      gt3_rxcharisk_out,
        gt3_rxdisperr_out               =>      gt3_rxdisperr_out,
        gt3_rxnotintable_out            =>      gt3_rxnotintable_out,
    ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt3_gtprxn_in                   =>      XAUI_RX_L3_N,
        gt3_gtprxp_in                   =>      XAUI_RX_L3_P,
    ------------------ Receive Ports - RX Channel Bonding Ports ----------------
        gt3_rxchanbondseq_out           =>      gt3_rxchanbondseq_out,
        gt3_rxchbonden_in               =>      '1',
        gt3_rxchbondi_in                =>      gt0_rxchbondo_out,
        gt3_rxchbondlevel_in            =>      "000",	-- no more daisy chaining
        gt3_rxchbondmaster_in           =>      '0',
        gt3_rxchbondo_out               =>      open,
        gt3_rxchbondslave_in            =>      '1',	-- 0 master, 1,2,3 slave
    ----------------- Receive Ports - RX Channel Bonding Ports  ----------------
        gt3_rxchanisaligned_out         =>      gt3_rxchanisaligned_out,
        gt3_rxchanrealign_out           =>      open,
    ------------ Receive Ports - RX Decision Feedback Equalizer(DFE) -----------
        gt3_dmonitorout_out             =>      open,
    -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt3_rxlpmhfhold_in              =>      '0',
        gt3_rxlpmhfovrden_in            =>      '0',
        gt3_rxlpmlfhold_in              =>      '0',
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt3_rxoutclkfabric_out          =>      open,
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt3_gtrxreset_in                =>      SYNC_RESET_CLK156,
        gt3_rxlpmreset_in               =>      '0',
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt3_rxpolarity_in               =>      gt_rxpolarity_in,
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt3_rxresetdone_out             =>      open,
    --------------------- TX Initialization and Reset Ports --------------------
        gt3_gttxreset_in                =>      SYNC_RESET_CLK156,
        gt3_txuserrdy_in                =>      GT_TXUSERRDY,
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt3_txdata_in                   =>      gt3_txdata_in,
    ------------------ Transmit Ports - TX 8B/10B Encoder Ports ----------------
        gt3_txcharisk_in                =>      gt3_txcharisk_in,
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
        gt3_gtptxn_out                  =>      XAUI_TX_L3_N,
        gt3_gtptxp_out                  =>      XAUI_TX_L3_P,
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt3_txoutclkfabric_out          =>      open,
        gt3_txoutclkpcs_out             =>      open,
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt3_txresetdone_out             =>      open,
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt3_txpolarity_in               =>      gt_txpolarity_in,

    --____________________________COMMON PORTS________________________________
   GT0_PLL0RESET_OUT  => GT0_PLL0RESET_OUT,
         GT0_PLL0OUTCLK_OUT  => open,
         GT0_PLL0OUTREFCLK_OUT  => open,
         GT0_PLL0LOCK_OUT  => CLK156_LOCK,
         GT0_PLL0REFCLKLOST_OUT  => open,
         GT0_PLL1OUTCLK_OUT  => open,
         GT0_PLL1OUTREFCLK_OUT  => open,
     sysclk_in => CLK156g	-- 10 MHz reference clock. Change XAUI core configuration from the default 100 MHz to 156.25 MHz

);
BUFG_003: BUFG  port map (I=> CLK156, O=> CLK156g);

XAUI_DEBUG(5) <= gt1_rxchanisaligned_out and gt2_rxchanisaligned_out and gt3_rxchanisaligned_out;
	-- bit5: FPGA XAUI receiver is synchronized across all 4 lanes (3 slaves aligned with 1 master)

gt_rxpolarity_in <= '0';	-- '0' no inversion, '1' inverted
gt_txpolarity_in <= '0';	-- '0' no inversion, '1' inverted




--//-- XGMII INTERFACE ---------------------------------
-- internal 64-bit wide SDR XGMII data path to/from the 10G Ethernet MAC.
-- mapping of lane to XGMII data bits

-- Byte order is 0,1,2,3,0,1,2,3
XAUI_RXD(7 downto 0) <= gt0_rxdata_out(7 downto 0);
XAUI_RXD(15 downto 8) <= gt1_rxdata_out(7 downto 0);
XAUI_RXD(23 downto 16) <= gt2_rxdata_out(7 downto 0);
XAUI_RXD(31 downto 24) <= gt3_rxdata_out(7 downto 0);
XAUI_RXD(39 downto 32) <= gt0_rxdata_out(15 downto 8);
XAUI_RXD(47 downto 40) <= gt1_rxdata_out(15 downto 8);
XAUI_RXD(55 downto 48) <= gt2_rxdata_out(15 downto 8);
XAUI_RXD(63 downto 56) <= gt3_rxdata_out(15 downto 8);

XAUI_RXCHARISK(3 downto 0) <= gt3_rxcharisk_out(0) & gt2_rxcharisk_out(0) & gt1_rxcharisk_out(0) & gt0_rxcharisk_out(0);
XAUI_RXCHARISK(7 downto 4) <= gt3_rxcharisk_out(1) & gt2_rxcharisk_out(1) & gt1_rxcharisk_out(1) & gt0_rxcharisk_out(1);
XAUI_RXDISPERR(3 downto 0) <= gt3_rxdisperr_out(0) & gt2_rxdisperr_out(0) & gt1_rxdisperr_out(0) & gt0_rxdisperr_out(0);
XAUI_RXDISPERR(7 downto 4) <= gt3_rxdisperr_out(1) & gt2_rxdisperr_out(1) & gt1_rxdisperr_out(1) & gt0_rxdisperr_out(1);
XAUI_RXNOTINTABLE(3 downto 0) <= gt3_rxnotintable_out(0) & gt2_rxnotintable_out(0) & gt1_rxnotintable_out(0) & gt0_rxnotintable_out(0);
XAUI_RXNOTINTABLE(7 downto 4) <= gt3_rxnotintable_out(1) & gt2_rxnotintable_out(1) & gt1_rxnotintable_out(1) & gt0_rxnotintable_out(1);

XAUI2XGMII_001: XAUI2XGMII PORT MAP(
	CLK => CLK156g,
	SYNC_RESET => SYNC_RESET_CLK156,
	XAUI_RXD => XAUI_RXD(31 downto 0),
	XAUI_RXCHARISK => XAUI_RXCHARISK(3 downto 0),
	XAUI_RXDISPERR => XAUI_RXDISPERR(3 downto 0),
	XAUI_RXNOTINTABLE => XAUI_RXNOTINTABLE(3 downto 0),
	XGMII_RXD => XGMII_RXD1(31 downto 0),
	XGMII_RXC => XGMII_RXC1(3 downto 0)
);

XAUI2XGMII_002: XAUI2XGMII PORT MAP(
	CLK => CLK156g,
	SYNC_RESET => SYNC_RESET_CLK156,
	XAUI_RXD => XAUI_RXD(63 downto 32),
	XAUI_RXCHARISK => XAUI_RXCHARISK(7 downto 4),
	XAUI_RXDISPERR => XAUI_RXDISPERR(7 downto 4),
	XAUI_RXNOTINTABLE => XAUI_RXNOTINTABLE(7 downto 4),
	XGMII_RXD => XGMII_RXD1(63 downto 32),
	XGMII_RXC => XGMII_RXC1(7 downto 4)
);

-- XGMII loopback
XGMII_RXD <= XGMII_RXD1 when (CREG(1)(0) = '0') else XGMII_TXD;
XGMII_RXC <= XGMII_RXC1 when (CREG(1)(0) = '0') else XGMII_TXC;


XGMII2XAUI_001: XGMII2XAUI
GENERIC MAP(
	NBYTES => 8
)
PORT MAP(
	CLK => CLK156g,
	SYNC_RESET => SYNC_RESET_CLK156,
	XGMII_TXD => XGMII_TXD,
	XGMII_TXC => XGMII_TXC,
	XAUI_TXD => XAUI_TXD,
	XAUI_TXCHARISK => XAUI_TXCHARISK
);

-- Byte order is 0,1,2,3,0,1,2,3
gt0_txdata_in(7 downto 0) <= XAUI_TXD(7 downto 0);
gt1_txdata_in(7 downto 0) <= XAUI_TXD(15 downto 8);
gt2_txdata_in(7 downto 0) <= XAUI_TXD(23 downto 16);
gt3_txdata_in(7 downto 0) <= XAUI_TXD(31 downto 24);
gt0_txdata_in(15 downto 8) <= XAUI_TXD(39 downto 32);
gt1_txdata_in(15 downto 8) <= XAUI_TXD(47 downto 40);
gt2_txdata_in(15 downto 8) <= XAUI_TXD(55 downto 48);
gt3_txdata_in(15 downto 8) <= XAUI_TXD(63 downto 56);

gt0_txcharisk_in <= XAUI_TXCHARISK(4) & XAUI_TXCHARISK(0);
gt1_txcharisk_in <= XAUI_TXCHARISK(5) & XAUI_TXCHARISK(1);
gt2_txcharisk_in <= XAUI_TXCHARISK(6) & XAUI_TXCHARISK(2);
gt3_txcharisk_in <= XAUI_TXCHARISK(7) & XAUI_TXCHARISK(3);

--//-- EXTERNAL PHY INTERFACE ---------------------------------
LEFT_CONNECTOR_A(1) <= LAN1_MDC;
LEFT_CONNECTOR_A(2) <= LAN1_MDIO_OUT when (LAN1_MDIO_DIR = '0') else 'Z';
LAN1_MDIO_IN <= LEFT_CONNECTOR_A(2);


-- PHY status monitoring  (must reclock otherwise Vivado's confused?)
MONITORING_001: process(CLK156g)
begin
	if rising_edge(CLK156g) then
		SREG(10)(0) <= not LEFT_CONNECTOR_A(4);	-- LASI
		SREG(10)(1) <= not LEFT_CONNECTOR_A(5);	-- RX link/activity
		SREG(10)(2) <= not LEFT_CONNECTOR_A(6);	-- TX link/activity
		SREG(10)(3) <= not LEFT_CONNECTOR_A(7);	-- SFP+ALARM
		SREG(10)(4) <= LEFT_CONNECTOR_A(8);	-- PGOOD 1.2V
		SREG(10)(5) <= LEFT_CONNECTOR_A(9);	-- PGOOD 3.3V
	end if;
end process;
LEFT_CONNECTOR_A(9 downto 4) <= (others => 'Z');

--//-- ETHERNET MAC#1  -----------------------------------
LAN1_MAC_ADDR_GEN: process(CLK156g)
begin
	if rising_edge(CLK156g) then
		LAN1_TEST_MODE(0) <= CREG(1)(1);	-- local loopback at the PHY
		--LAN1_TEST_MODE(1) <= CREG(1)(2);	future REMOTE LOOPBACK
		LAN1_PHY_RESET <= CREG(1)(6);	-- PHY soft reset
		LAN1_POWER_DOWN <= CREG(1)(4);	-- PHY power down

		-- MAC address automatically generated from unique DNA_ID
		if(DNA_ID_SAMPLE_CLK = '1') then
			LAN1_MAC_ADDR <= x"00" & DNA_ID_DATA(39 downto 0);	-- unique, unicast
		end if;
	end if;
end process;

-- simulate tx frame
LAN1_MAC_TX_SIM_001: if(SIMULATION = '1') generate
SIM_001: process(CLK156g)
begin
	if rising_edge(CLK156g) then
		TEST_CLK_CNTR <= TEST_CLK_CNTR + 1;
		case(to_integer(TEST_CLK_CNTR)) is
			when 14080 =>
				LAN1_MAC_TX_DATA <= x"0706050403020100";
				LAN1_MAC_TX_DATA_VALID <= x"FF";
			when 14081 =>
				LAN1_MAC_TX_DATA <= x"1716151413121110";
				LAN1_MAC_TX_DATA_VALID <= x"FF";
				LAN1_MAC_TX_EOF <= '1';
			when others =>
				LAN1_MAC_TX_DATA <= x"0000000000000000";
				LAN1_MAC_TX_DATA_VALID <= x"00";
				LAN1_MAC_TX_EOF <= '0';
		end case;
	end if;
end process;
end generate;

-- send a test Ethernet frame once per second
LAN1_MAC_TX_001: if(SIMULATION = '0') generate
TEST_001: process(CLK156g)
begin
	if rising_edge(CLK156g) then
		TICK_1S_SHIFT(0) <= TICK_1S;
		TICK_1S_SHIFT(6 downto 1) <= TICK_1S_SHIFT(5 downto 0);

		if(TICK_1S = '1') then
			-- Byte order: LSB first
			LAN1_MAC_TX_DATA <= x"0E00FFFFFFFFFFFF";	-- preamble + broadcast address + source address
			LAN1_MAC_TX_DATA_VALID <= x"FF";
			LAN1_MAC_TX_EOF <= '0';
		elsif(TICK_1S_SHIFT(0) = '1') then
			LAN1_MAC_TX_DATA <= x"01000608A3BBCA08";	-- source address
		elsif(TICK_1S_SHIFT(1) = '1') then
			LAN1_MAC_TX_DATA <= x"0E00010004060008";	-- data
		elsif(TICK_1S_SHIFT(2) = '1') then
			LAN1_MAC_TX_DATA <= x"7E0110ACA3BBCA08";	-- data
		elsif(TICK_1S_SHIFT(3) = '1') then
			LAN1_MAC_TX_DATA <= x"10AC000000000000";	-- data
		elsif(TICK_1S_SHIFT(4) = '1') then
			LAN1_MAC_TX_DATA <= x"0000000000001F01";	-- data
-- TEST TEST TEST
			LAN1_MAC_TX_DATA_VALID <= x"03";
			LAN1_MAC_TX_EOF <= '1';

--		elsif(TICK_1S_SHIFT(5) = '1') then
--			LAN1_MAC_TX_DATA <= x"0000000000000000";	-- data
--		elsif(TICK_1S_SHIFT(6) = '1') then
--			LAN1_MAC_TX_DATA <= x"D3C41B1300000000";	-- data
--			LAN1_MAC_TX_EOF <= '1';
		else
			LAN1_MAC_TX_DATA <= (others => '0');
			LAN1_MAC_TX_DATA_VALID <= (others => '0');
			LAN1_MAC_TX_EOF <= '0';
		end if;
	end if;
end process;
end generate;


COM5501_001: COM5501
GENERIC MAP(
	EXT_PHY_MDIO_ADDR => "00000",	-- on COM-5104 adapter, the external PHY MDIO address is 0
	RX_MTU => 1500,	-- bytes in standard frame
	RX_BUFFER => '1',	-- minimize latency. No rx output buffer, use same clock for CLK and CLK156g.
	RX_BUFFER_ADDR_NBITS => 10,	-- n/a
	TX_MTU => 1500,	-- bytes in standard frame
	TX_BUFFER => '1',	-- minimize latency. No tx input buffer, use same clock for CLK and CLK156g.
	TX_BUFFER_ADDR_NBITS => 10,	-- n/a
	MAC_CONTROL_PAUSE_ENABLE => '1',
	SIMULATION => SIMULATION
)
PORT MAP(
	CLK => CLK156g,
		-- In this example we use the same 156.25 MHz clock as user clock,
		-- it does not have to be so.
	SYNC_RESET => SYNC_RESET_CLK156,
	CLK156g => CLK156g,
	MAC_TX_CONFIG => x"03",	-- short frame padding,
	MAC_RX_CONFIG => x"0F",
	MAC_ADDR => LAN1_MAC_ADDR,
	MAC_TX_DATA => LAN1_MAC_TX_DATA,
	MAC_TX_DATA_VALID => LAN1_MAC_TX_DATA_VALID,
	MAC_TX_EOF => LAN1_MAC_TX_EOF,
	MAC_TX_CTS => LAN1_MAC_TX_CTS,
	MAC_RX_DATA => open,
	MAC_RX_DATA_VALID => open,
	MAC_RX_SOF => open,
	MAC_RX_EOF => open,
	MAC_RX_FRAME_VALID => open,
	MAC_RX_CTS => '1',
	-- XGMII interface
	XGMII_TXD => XGMII_TXD,
	XGMII_TXC => XGMII_TXC,
	XGMII_RXD => XGMII_RXD,
	XGMII_RXC => XGMII_RXC,
	-- MDIO interface with external PHY
	RESET_N => LEFT_CONNECTOR_A(3),	-- pulse must be > 100ns (VSC8486-11)
	MDC => LAN1_MDC,
	MDIO_OUT => LAN1_MDIO_OUT,
	MDIO_IN => LAN1_MDIO_IN,
	MDIO_DIR => LAN1_MDIO_DIR,
	PHY_CONFIG_CHANGE => PHY_CONFIG_CHANGE,	-- MANDATORY in many cases (for example when inverted differential traces)
	PHY_RESET => LAN1_PHY_RESET,
	TEST_MODE => LAN1_TEST_MODE,
	POWER_DOWN => LAN1_POWER_DOWN,
	PHY_STATUS => LAN1_PHY_STATUS,
	PHY_STATUS2 => LAN1_PHY_STATUS2,
	PHY_ID => LAN1_PHY_ID,
	N_TX_FRAMES => LAN1_N_TX_FRAMES,
	N_RX_FRAMES => LAN1_N_RX_FRAMES,
	N_RX_BAD_CRCS => LAN1_N_RX_BAD_CRCS,
	N_RX_FRAMES_TOO_SHORT => open,
	N_RX_FRAMES_TOO_LONG => open,
	N_RX_WRONG_ADDR => open,
	N_RX_LENGTH_ERRORS => open,
	RX_IPG => LAN1_RX_IPG,
	DEBUG1 => DEBUG1,
	DEBUG2 => DEBUG2,
	DEBUG3 => DEBUG3,
	TP => LAN1_TP
);
PHY_CONFIG_CHANGE <= CONFIG_CHANGE_PULSE;

-- PHY status monitoring
MONITORING_002: process(CLK156g)
begin
	if rising_edge(CLK156g) then
		SREG(11) <= LAN1_PHY_ID(7 downto 0);	-- PHY device ID. Expecting 0x8486 with VSC8486-11
		SREG(12) <= LAN1_PHY_ID(15 downto 8);	-- PHY device ID. Expecting 0x8486 with VSC8486-11
		SREG(13) <= LAN1_PHY_STATUS2;	-- PHY SFP+ side status.
		SREG(14) <= LAN1_PHY_STATUS;	-- PHY XAUI rx status. Expecting 0x3F
			-- bit0: all PHY XAUI rx lanes in sync
			-- bit1: PHY XAUI rx PLL in lock
			-- bit2: PHY XAUI rx lane0 signal present
			-- bit3: PHY XAUI rx lane1 signal present
			-- bit4: PHY XAUI rx lane2 signal present
			-- bit5: PHY XAUI rx lane3 signal present
		SREG(15)(5 downto 0) <= XAUI_DEBUG;	-- FPGA XAUI status.
			-- bit5: FPGA XAUI receiver is synchronized across all 4 lanes
		--SREG(16) <= ;
            -- bit 0:
		SREG(17) <= LAN1_N_RX_FRAMES(7 downto 0);
		SREG(18) <= LAN1_N_RX_FRAMES(15 downto 8);
		SREG(19) <= LAN1_N_RX_BAD_CRCS(7 downto 0);
		SREG(20) <= LAN1_N_RX_BAD_CRCS(15 downto 8);
		SREG(21) <= LAN1_RX_IPG;

		SREG(22) <= LAN1_MAC_ADDR(47 downto 40);
		SREG(23) <= LAN1_MAC_ADDR(39 downto 32);
		SREG(24) <= LAN1_MAC_ADDR(31 downto 24);
		SREG(25) <= LAN1_MAC_ADDR(23 downto 16);
		SREG(26) <= LAN1_MAC_ADDR(15 downto 8);
		SREG(27) <= LAN1_MAC_ADDR(7 downto 0);
			-- local MAC address

--		if(LATCH_MONITORING_PULSE = '1') then
			SREG(28) <= DEBUG1(7 downto 0);
			SREG(29) <= DEBUG1(15 downto 8);
			SREG(30) <= DEBUG1(23 downto 16);
			SREG(31) <= DEBUG1(31 downto 24);
			SREG(32) <= DEBUG1(39 downto 32);
			SREG(33) <= DEBUG1(47 downto 40);
			SREG(34) <= DEBUG1(55 downto 48);
			SREG(35) <= DEBUG1(63 downto 56);

			SREG(36) <= DEBUG2(7 downto 0);
			SREG(37) <= DEBUG2(15 downto 8);
			SREG(38) <= DEBUG2(23 downto 16);
			SREG(39) <= DEBUG2(31 downto 24);
			SREG(40) <= DEBUG2(39 downto 32);
			SREG(41) <= DEBUG2(47 downto 40);
			SREG(42) <= DEBUG2(55 downto 48);
			SREG(43) <= DEBUG2(63 downto 56);

			SREG(44) <= DEBUG3(7 downto 0);
			SREG(45) <= DEBUG3(15 downto 8);
			SREG(46) <= DEBUG3(23 downto 16);
			SREG(47) <= DEBUG3(31 downto 24);
			SREG(48) <= DEBUG3(39 downto 32);
			SREG(49) <= DEBUG3(47 downto 40);
			SREG(50) <= DEBUG3(55 downto 48);
			SREG(51) <= DEBUG3(63 downto 56);
--		end if;
	end if;
end process;


RX_LAN_BUFFER_EMPTY <= '1'; -- until 10G MAC code in place


--// TEST POINTS  -----------------------------------------------
-- Warning: test points can make timing much worse!
RIGHT_CONNECTOR_A(10 downto 1) <= LAN1_TP;
RIGHT_CONNECTOR_A(16 downto 11) <= XAUI_DEBUG(5 downto 0);
RIGHT_CONNECTOR_A(17) <= CONFIG_CHANGE_PULSE;


--// ARM CO-PROCESSOR INTERFACE ---------------------------------------------------
-- Primarily used for monitoring and control.
-- 8-bit shared address/data bus. clock synchronous.
-- PART OF THE FRAMEWORK. DO NOT CHANGE unless you want to add more control registers
--(see UC_WRITE_001) or status registers (see UC_READ_001).
--
-- Address latch
UC_ADDR_001: process(UC_CSIB_IN, UC_WEBG, UC_ALE_IN, UC_AD)
begin
	if rising_edge(UC_WEBG) then
		if (UC_CSIB_IN = '0') and (UC_ALE_IN = '1') then
			UC_ADDRESS <= unsigned(UC_AD);
	  	end if;
  	end if;
end process;

-- Read status registers
-- User can define additional control registers using the same pattern.
UC_READ_001: process(UC_ADDRESS, REG255, RX_LAN, SREG)
begin
	case(UC_ADDRESS) is
		-- ComBlock-reserved addresses ----
		when "11111111" => UC_AD_LOCAL <= REG255;		-- reg 255. Async serial from 3 connectors
		when "11111110" => UC_AD_LOCAL <= RX_LAN;-- reg 254 = 8-bit data from LAN M&C channel
		when "11111101" => UC_AD_LOCAL <= REVISION;	-- reg 253 = fpga revision
		when "11111100" => UC_AD_LOCAL <= OPTION;		-- reg 252 = fpga option

		-- User-defined status registers -------
		-- SREG0-6 reserved for use by the ARM microcontroller
		when "00000111" => UC_AD_LOCAL <= SREG(7);
		when "00001000" => UC_AD_LOCAL <= SREG(8);
		when "00001001" => UC_AD_LOCAL <= SREG(9);
		when "00001010" => UC_AD_LOCAL <= SREG(10);
		when "00001011" => UC_AD_LOCAL <= SREG(11);
		when "00001100" => UC_AD_LOCAL <= SREG(12);
		when "00001101" => UC_AD_LOCAL <= SREG(13);
		when "00001110" => UC_AD_LOCAL <= SREG(14);
		when "00001111" => UC_AD_LOCAL <= SREG(15);
		when "00010000" => UC_AD_LOCAL <= SREG(16);
		when "00010001" => UC_AD_LOCAL <= SREG(17);
		when "00010010" => UC_AD_LOCAL <= SREG(18);
		when "00010011" => UC_AD_LOCAL <= SREG(19);
		when "00010100" => UC_AD_LOCAL <= SREG(20);
		when "00010101" => UC_AD_LOCAL <= SREG(21);
		when "00010110" => UC_AD_LOCAL <= SREG(22);
		when "00010111" => UC_AD_LOCAL <= SREG(23);
		when "00011000" => UC_AD_LOCAL <= SREG(24);
		when "00011001" => UC_AD_LOCAL <= SREG(25);
		when "00011010" => UC_AD_LOCAL <= SREG(26);
		when "00011011" => UC_AD_LOCAL <= SREG(27);
		when "00011100" => UC_AD_LOCAL <= SREG(28);
		when "00011101" => UC_AD_LOCAL <= SREG(29);
		when "00011110" => UC_AD_LOCAL <= SREG(30);
		when "00011111" => UC_AD_LOCAL <= SREG(31);
		when "00100000" => UC_AD_LOCAL <= SREG(32);
		when "00100001" => UC_AD_LOCAL <= SREG(33);
		when "00100010" => UC_AD_LOCAL <= SREG(34);
		when "00100011" => UC_AD_LOCAL <= SREG(35);
		when "00100100" => UC_AD_LOCAL <= SREG(36);
		when "00100101" => UC_AD_LOCAL <= SREG(37);
		when "00100110" => UC_AD_LOCAL <= SREG(38);
		when "00100111" => UC_AD_LOCAL <= SREG(39);
		when "00101000" => UC_AD_LOCAL <= SREG(40);
		when "00101001" => UC_AD_LOCAL <= SREG(41);
		when "00101010" => UC_AD_LOCAL <= SREG(42);
		when "00101011" => UC_AD_LOCAL <= SREG(43);
		when "00101100" => UC_AD_LOCAL <= SREG(44);
		when "00101101" => UC_AD_LOCAL <= SREG(45);
		when "00101110" => UC_AD_LOCAL <= SREG(46);
		when "00101111" => UC_AD_LOCAL <= SREG(47);
		when "00110000" => UC_AD_LOCAL <= SREG(48);
		when "00110001" => UC_AD_LOCAL <= SREG(49);
		when "00110010" => UC_AD_LOCAL <= SREG(50);
		when "00110011" => UC_AD_LOCAL <= SREG(51);


		-- user can add more status registers as needed (200+)
		when others => UC_AD_LOCAL <= (others => '0');
	end case;
end process;

UC_AD <= UC_AD_LOCAL when (UC_CSIB_IN = '0') and (UC_REB_IN = '0') else (others => 'Z');
	-- when to drive the data bus between ARM and FPGA

-- toggle a few flags upon reading specific status registers
UC_READ_002: process(ASYNC_RESET, UC_REBG, UC_CSIB_IN, UC_ADDRESS,
						SREG254_READ_TOGGLE)
begin
	if(ASYNC_RESET = '1') then
		SREG254_READ_TOGGLE <= '0';
	elsif rising_edge(UC_REBG) then
		if (UC_CSIB_IN = '0')  then
			if (UC_ADDRESS = 7) then
				SREG7_READ_TOGGLE <= not SREG7_READ_TOGGLE;
			end if;
			if (UC_ADDRESS = 254) then
				SREG254_READ_TOGGLE <= not SREG254_READ_TOGGLE;
			end if;
		end if;
	end if;
end process;

-- reclock with CLK156g
RECLOCK_SREG9_TOGGLE: process(CLK156g,SREG7_READ_TOGGLE)
begin
	if rising_edge(CLK156g) then
		SREG7_READ_TOGGLE_D <= SREG7_READ_TOGGLE;
		SREG7_READ_TOGGLE_D2 <= SREG7_READ_TOGGLE_D;
		if(SREG7_READ_TOGGLE_D /= SREG7_READ_TOGGLE_D2) then
			LATCH_MONITORING_PULSE <= '1';
		else
			LATCH_MONITORING_PULSE <= '0';
		end if;
	end if;
end process;

-- write to FPGA control registers
-- Users can define control registers as needed (up to 230) by modifying the UC_WRITE_001 process below.
UC_WRITE_001ax: if (SIMULATION = '0') generate
	UC_WRITE_001a: process(UC_WEBG)
	begin
		if rising_edge(UC_WEBG) then
			if (UC_CSIB_IN = '0') and (UC_ALE_IN = '0') and (UC_REB_IN = '1')  then
				for I in NCREG_IMIN to NCREG_IMAX loop
					if(UC_ADDRESS = I) then
						CREG(I) <= UC_AD;
					end if;
				end loop;
			end if;
		end if;
	end process;

	UC_WRITE_001: process(UC_CSIB_IN, UC_WEBG, UC_ALE_IN, UC_REB_IN, UC_AD)
	begin
		if rising_edge(UC_WEBG) then
			if (UC_CSIB_IN = '0') and (UC_ALE_IN = '0') and (UC_REB_IN = '1')  then

				if (UC_ADDRESS = NCREG_IMAX) then
					-- dummy write to last control register
					CONFIG_CHANGE_TOGGLE <= not CONFIG_CHANGE_TOGGLE;
					-- Configuration change toggles upon writing the last control register
					-- This happens invisibly to the user (only the ARM uC writes to this last control register
					-- which is invible to the user and to the ComBlock Control Center).
				end if;

				-- Reserved:
				-- REG254 reserved for output serial
				-- REG255 write reserved for output serial (8-bit parallel format)
			end if;
		end if;
	end process;
end generate;


-- initialize control registers for simulation. Ignored at runtime.
UC_WRITE_001y: if (SIMULATION = '1') generate
process
begin
	CREG(0) <= x"00";
	CREG(1) <= x"00";
	CREG(2) <= x"00";
	CREG(3) <= x"00";
	CREG(4) <= x"00";
	CREG(5) <= x"00";
	CREG(6) <= x"01";
	CREG(7) <= x"00";
	CONFIG_CHANGE_TOGGLE <= '0';
	-- etc
	wait for 66us;
	CONFIG_CHANGE_TOGGLE <= '1';
	wait for 134us;
	CONFIG_CHANGE_TOGGLE <= '0';

	wait;
end process;

end generate;

-- Reclock CONFIG_CHANGE_TOGGLE to be synchronous with processing clock CLK156g
RECLOCK_002: process(CLK156g)
begin
	if rising_edge(CLK156g) then
		CONFIG_CHANGE_TOGGLE_D <= CONFIG_CHANGE_TOGGLE;
		CONFIG_CHANGE_TOGGLE_D2 <= CONFIG_CHANGE_TOGGLE_D;
		if(CONFIG_CHANGE_TOGGLE_D /= CONFIG_CHANGE_TOGGLE_D2) then
			CONFIG_CHANGE_PULSE <= '1';
		else
			CONFIG_CHANGE_PULSE <= '0';
		end if;
	end if;
end process;

-- DNA Port ------------------------------------
-- Read FPGA unique DNA ID
DNA_ID_001: DNA_ID
	GENERIC MAP(
		CLK_FREQUENCY => CLK_FREQUENCY	-- CLK156g in MHz, as time reference
	)
	PORT MAP(
		CLK => CLK156g,
		SYNC_RESET => SYNC_RESET_CLK156,
		ID_OUT => DNA_ID_DATA,
		ID_VALID_OUT => open,
		ID_SAMPLE_CLK_OUT => DNA_ID_SAMPLE_CLK
);


-- M&C USB interface --------------------------
-- REG255 reserved for reading serial port inputs
-- These signals are pulled high (to mimic stop bit).
REG255 <= "1111" & RX_LAN_BUFFER_EMPTY & "111";
	-- M&C port through LAN
	-- indicates AVAILABILITY of 8-bit byte from LAN. Not actual data.
	-- When low, uC must read byte from LAN


-- Immediately upon completing reading a M&C byte from the USB or LAN, ask for the
-- next one.
RECLOCK_RDN_D: process(CLK156g, SREG254_READ_TOGGLE)
begin
	if rising_edge(CLK156g) then
		SREG254_READ_TOGGLE_D <= SREG254_READ_TOGGLE;
		SREG254_READ_TOGGLE_D2 <= SREG254_READ_TOGGLE_D;

		RX_LAN_BUFFER_EMPTY_D <= RX_LAN_BUFFER_EMPTY;
		RX_LAN_BUFFER_EMPTY_D2 <= RX_LAN_BUFFER_EMPTY_D;


		if (SREG254_READ_TOGGLE_D2 /= SREG254_READ_TOGGLE_D) then
			-- end of M&C byte read from ARM uC.
			if(RX_LAN_BUFFER_EMPTY_D2 = '0') then
				-- last M&C byte read was over LAN. Increment LAN elastic buffer read pointer
				RX_LAN_SAMPLE_CLK_REQ <= '1';
					-- identifies LAN as the media through which	this module exchanges
					-- M&C information. Response will be directed the same way.
			end if;
		else
			RX_LAN_SAMPLE_CLK_REQ <= '0';
		end if;
	end if;
end process;

end Behavioral;
